//
// FX68K
//
// M68K cycle accurate, fully synchronous
// Copyright 2018 by Jorge Cwik
//
module nanoRom( input clk, input [9-1:0] nanoAddr, output reg [68-1:0] nanoOutput);

  always @( posedge clk)
  begin
    case (nanoAddr)
      9'h  0: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h  1: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h  2: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h  3: nanoOutput = 68'b00000000000000000000000000001000000110011100000000000000101001000001;
      9'h  4: nanoOutput = 68'b00100001000000011000010001001000000110100000000001000000011001001001;
      9'h  5: nanoOutput = 68'b00000001100000000010100000001000000110000000001001000000001001001001;
      9'h  6: nanoOutput = 68'b00100000000000011000010001000000000101000000000010000000100001010000;
      9'h  7: nanoOutput = 68'b11000001000000000000000000001000000100010000000001000000000001010001;
      9'h  8: nanoOutput = 68'b00100001000000011000010000000000000000000000000101000000000000010000;
      9'h  9: nanoOutput = 68'b01000001011000000000100000000110010001000000001100000000110100011000;
      9'h  a: nanoOutput = 68'b01000001011000000000100000000110010001000000001100000001100100011000;
      9'h  b: nanoOutput = 68'b00100001000000011000010000000000000100000000000001000000000001010000;
      9'h  c: nanoOutput = 68'b10100100001000011000001000010000101001110000000001000100110010100001;
      9'h  d: nanoOutput = 68'b01000000000000000000000010000000010100000000001000110001000000000000;
      9'h  e: nanoOutput = 68'b00100001000000011000000000110010100100011111010001100000000001000000;
      9'h  f: nanoOutput = 68'b00100010000000011000000000000000100010000100000000010100000100000011;
      9'h 10: nanoOutput = 68'b00000001011000000000000001000110000000000000000010000000000100000000;
      9'h 11: nanoOutput = 68'b00000000000000000000000000001000000100000000000001000000000001010001;
      9'h 12: nanoOutput = 68'b00000001100000000010100000001000000110000000001001010000001001001001;
      9'h 13: nanoOutput = 68'b00101000000000001000010000000000000000000000000010000000000000000000;
      9'h 14: nanoOutput = 68'b01100010000000011000010010000000010100000000001000110001000000000000;
      9'h 15: nanoOutput = 68'b00000000000000000000000010010010100000000000000100110010000000000000;
      9'h 16: nanoOutput = 68'b00100000000000011000010001001000000110000000001001010000001001001001;
      9'h 17: nanoOutput = 68'b00000000000000000000001000000000100100000000000000110010000001011000;
      9'h 18: nanoOutput = 68'b00010010000000000100100000001000000100000000000010000000000001010001;
      9'h 19: nanoOutput = 68'b00100010000000011100000000000000000001100000000010001000100000000000;
      9'h 1a: nanoOutput = 68'b00010010000000000100000000000000010001100000000010000000000000000000;
      9'h 1b: nanoOutput = 68'b00000000000000000000000000011001100110100000010001000000011011010001;
      9'h 1c: nanoOutput = 68'b10100010110000000000000000000000100000010000010010000100000100000000;
      9'h 1d: nanoOutput = 68'b10000000000000000000000000001000000100010000000001000000000001000001;
      9'h 1e: nanoOutput = 68'b00100000000000011001000000011010000110000000001001000000001001001001;
      9'h 1f: nanoOutput = 68'b00010011000000000000101000010000001001000000010101000000100000110000;
      9'h 20: nanoOutput = 68'b00000001000000000001010000000000000000000000000101100000000000010000;
      9'h 21: nanoOutput = 68'b00100010000000011000001000001000100110000000000001000000000001010001;
      9'h 22: nanoOutput = 68'b00000001000000000010100001010000001001000000010110000000100000110000;
      9'h 23: nanoOutput = 68'b01000001000000000000000000000000000001101010001100000000110000000000;
      9'h 24: nanoOutput = 68'b00110100000000000100000100000000000000000000000010000000000000000000;
      9'h 25: nanoOutput = 68'b00000000000100100000100000000000010000000000000000000001000000011000;
      9'h 26: nanoOutput = 68'b01110101000000000100100000100010000001100000000000000000110100001010;
      9'h 27: nanoOutput = 68'b00100010000000011010000100000000100010000100000000010100000100000011;
      9'h 28: nanoOutput = 68'b11000001000000000000000000001000000100010000000001000000000001010001;
      9'h 29: nanoOutput = 68'b01010011000000000100100000100010000001100000000000000000110100001010;
      9'h 2a: nanoOutput = 68'b11000001000000000000000000001001100110110000000001000000011011000001;
      9'h 2b: nanoOutput = 68'b01001001110000000000001000001000001000000000000101000000000000100001;
      9'h 2c: nanoOutput = 68'b00000000000000000000100000100010010000000000000000110001000100000010;
      9'h 2d: nanoOutput = 68'b00010000110000000001010000000000000000011100000010000000000000011000;
      9'h 2e: nanoOutput = 68'b01010001110000000001000000011010100100000000000001000000000001000001;
      9'h 2f: nanoOutput = 68'b00000000000000000000000001000000000100000000001100010000000001010000;
      9'h 30: nanoOutput = 68'b00001000000000011001001000001000000110100000000001000100000011010001;
      9'h 31: nanoOutput = 68'b01010001110000000001010000001000001000000000000101000000000000110001;
      9'h 32: nanoOutput = 68'b10100010110100100100000001000000000001110000000010000000110000010000;
      9'h 33: nanoOutput = 68'b00000000000100000000000000000010100001001010000101100000100000010000;
      9'h 34: nanoOutput = 68'b00010000110000000001000000000000100000000000010010000100000100000000;
      9'h 35: nanoOutput = 68'b10000000000000000000000000001000000100010000000001000000000001000001;
      9'h 36: nanoOutput = 68'b00000001000000000000000001000000001001000000000101000000100000100000;
      9'h 37: nanoOutput = 68'b00010010000000000000100000001010101000000000000101000000000000110001;
      9'h 38: nanoOutput = 68'b10100000000100111000000000100001100010111010000101100000011010010010;
      9'h 39: nanoOutput = 68'b00100000000000011000000000110010100110000000010000100000001101000010;
      9'h 3a: nanoOutput = 68'b00010010000000001100000000000000000000000000000010000000000000000000;
      9'h 3b: nanoOutput = 68'b11000001000000000000001000011101100100010000000001000000000001000001;
      9'h 3c: nanoOutput = 68'b00010100000000000100000100000000000000000000000010000000000000000000;
      9'h 3d: nanoOutput = 68'b10100010110000000100001000000000100000010000010010000100000010000000;
      9'h 3e: nanoOutput = 68'b00100000000100111000000000000000100000010010000101000100000100010010;
      9'h 3f: nanoOutput = 68'b00100010000000011000000000000000100010000100000000010100000100000011;
      9'h 40: nanoOutput = 68'b00100010100000011001010000010000100100000000001110000100001000000000;
      9'h 41: nanoOutput = 68'b00000000000100000000000000000010100000001010000101000000000000010000;
      9'h 42: nanoOutput = 68'b00100010100000011001000000010010100100000000001110000100001000000000;
      9'h 43: nanoOutput = 68'b00000001000000000000010000000000100000000000010101000100000010010000;
      9'h 44: nanoOutput = 68'b00000000000100100000000000100010000000000100000000110001000100011010;
      9'h 45: nanoOutput = 68'b00100000000000011000000000010000100110000000011000100000001001000000;
      9'h 46: nanoOutput = 68'b00000000000100100000100000100010010000000000000000110001000100011010;
      9'h 47: nanoOutput = 68'b00000000011000000000000000000110000000000000001110000000110100111000;
      9'h 48: nanoOutput = 68'b00011000000000011001001000001000000100000000000001000000000001010001;
      9'h 49: nanoOutput = 68'b00100010000000011100000000000000000001100000000010001000100000000000;
      9'h 4a: nanoOutput = 68'b00110000100000001000000100000000100000000000000010000100000100000000;
      9'h 4b: nanoOutput = 68'b00000000000100000000000000000010100001000000000101100000100000010000;
      9'h 4c: nanoOutput = 68'b10100010110000000100001000010001100000010000000010000000000000000000;
      9'h 4d: nanoOutput = 68'b01000001000000000000000000000000000000000000000101000000000000010000;
      9'h 4e: nanoOutput = 68'b10000000000000000000000000001000000100010000000001000000000001000001;
      9'h 4f: nanoOutput = 68'b00000000000000000000000000001000001000000000000101000000000000110001;
      9'h 50: nanoOutput = 68'b00001000110000000000001000000000000000000000000010000000000000000000;
      9'h 51: nanoOutput = 68'b00010010000000001100000000000000000000000000000010000000000000000000;
      9'h 52: nanoOutput = 68'b00010000000000001010000100000000110001000000000010000100011000000000;
      9'h 53: nanoOutput = 68'b01010001000000011000001000000000000001100000000000000000110000000000;
      9'h 54: nanoOutput = 68'b00001100000000011000001000100001000010100000000101110000000000000011;
      9'h 55: nanoOutput = 68'b01000000000000000000000010000000010100000000001000110000000001000000;
      9'h 56: nanoOutput = 68'b11000001000000000000000000001000001000010000000101000000000000100001;
      9'h 57: nanoOutput = 68'b00000000000000000000000000001000000100011100000001100000000001000001;
      9'h 58: nanoOutput = 68'b00000000000000000000000000000000000000000000000101100000000000000000;
      9'h 59: nanoOutput = 68'b00000000000100000000000000000000100000000000000101000100000100010000;
      9'h 5a: nanoOutput = 68'b11101011000000000000000000000000000000010000000010000000000000000000;
      9'h 5b: nanoOutput = 68'b01100001000000011001000000011010100100000000000001000000000001000001;
      9'h 5c: nanoOutput = 68'b01100010000000011000010010000000010100000000001000110000000001000000;
      9'h 5d: nanoOutput = 68'b00000000000000000000000010010010100000000000010100110000000100000000;
      9'h 5e: nanoOutput = 68'b01000001000000000000010000011001101000000000000101000100001000110001;
      9'h 5f: nanoOutput = 68'b00100000000100111100000000000000000010000010000100100010001000010000;
      9'h 60: nanoOutput = 68'b00010010000000000000000000000010110100000000001110000000000000011000;
      9'h 61: nanoOutput = 68'b00000000000000000000001000010000100100000000011100110010000001011000;
      9'h 62: nanoOutput = 68'b00000000000100000000000000010000111000000000010101000100011000110000;
      9'h 63: nanoOutput = 68'b00000000011000000010100000000110000100000000001101110000000101000000;
      9'h 64: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h 65: nanoOutput = 68'b00000001000000000000000000000000010101001010001101000000100001010000;
      9'h 66: nanoOutput = 68'b00000001000000000000010000000000100000000000000101000100001000010000;
      9'h 67: nanoOutput = 68'b01110101000000010000001000000000000001100000000000000000110000000000;
      9'h 68: nanoOutput = 68'b01000001000000000000000010000000010100001010001000110001000000000000;
      9'h 69: nanoOutput = 68'b00100010000000011000000000011010101010000000010101000000001100110001;
      9'h 6a: nanoOutput = 68'b00100001000000011000010001010000000100000000010000010000000001010000;
      9'h 6b: nanoOutput = 68'b01000001000000000000010000000000100000000110000101000000000000010000;
      9'h 6c: nanoOutput = 68'b01000001000000000000000010000000010100001010001000110001000000000000;
      9'h 6d: nanoOutput = 68'b00100000000000011000010001010001000000000000011010000000000010001000;
      9'h 6e: nanoOutput = 68'b00000001000000000000000001010000000100000000010001110000000001000000;
      9'h 6f: nanoOutput = 68'b00010010000000001000000000011010101000000000000101000000000000110001;
      9'h 70: nanoOutput = 68'b00000000000000000000000000001000001000000000000101000000000000110001;
      9'h 71: nanoOutput = 68'b00010010000000000001100000000010000000000000000101100000000000000000;
      9'h 72: nanoOutput = 68'b00010010000000000001000000000010000100000000000101100000000000000000;
      9'h 73: nanoOutput = 68'b00100010000000011100000000001000001000000000000101000000000000100001;
      9'h 74: nanoOutput = 68'b00000001000000000001010000000000001010100000000110000000011000101000;
      9'h 75: nanoOutput = 68'b00000001100000000000100000000000000000000000000101000000000000010000;
      9'h 76: nanoOutput = 68'b00010010000000000000101000001001000100000000001001000000000011010001;
      9'h 77: nanoOutput = 68'b11110101001000000100000000000000000000010000000010000000000000000000;
      9'h 78: nanoOutput = 68'b00000000000000000000010000001001101000000000000101000010000010110001;
      9'h 79: nanoOutput = 68'b00000000000000000000010000000000100000000110000101100000000000000000;
      9'h 7a: nanoOutput = 68'b00100010100000001001100000000010000010000100001000000000001000001000;
      9'h 7b: nanoOutput = 68'b00100010100000001001000000000010000110000100001000000000001000001000;
      9'h 7c: nanoOutput = 68'b00010010000000001000010000000000000000000000001110000000000000011000;
      9'h 7d: nanoOutput = 68'b00110100000100101100000000000000000001100000000001100000110000010000;
      9'h 7e: nanoOutput = 68'b01110101000000001000000100000000111000000000010010000100000100000000;
      9'h 7f: nanoOutput = 68'b01000000000000000000010000010000100110000000011100100000000001011000;
      9'h 80: nanoOutput = 68'b11010011000000000000101000001001000100010000001001000000000011010001;
      9'h 81: nanoOutput = 68'b11110101001000000000000000000000100000010000000010000100000100000000;
      9'h 82: nanoOutput = 68'b01110101000000000100000000000000010000000000010010001000000001000000;
      9'h 83: nanoOutput = 68'b01110101000000000000000000000000110000000000010010001100000101000000;
      9'h 84: nanoOutput = 68'b01110101000000000000000000000000110000000000010010001100011001000000;
      9'h 85: nanoOutput = 68'b01110000000000011100000000000000000001100000001101000000110000000000;
      9'h 86: nanoOutput = 68'b00010000000000001000000000000010100000000000000010000000000000000000;
      9'h 87: nanoOutput = 68'b00010010000000000100000100000000010001000000000010000000000000000000;
      9'h 88: nanoOutput = 68'b01000000000000000000010000010000100110000000011100100010001001011000;
      9'h 89: nanoOutput = 68'b00100000000000011000010000000000000100000000000000100000000001000000;
      9'h 8a: nanoOutput = 68'b00000001000000000000000000000000001000000000000101000000000000110000;
      9'h 8b: nanoOutput = 68'b00100001000000011100000001011001000110000000011000000000001011001001;
      9'h 8c: nanoOutput = 68'b01100001000000011000000000010010100110000000011100100000001101011000;
      9'h 8d: nanoOutput = 68'b01100001000000011000010000010010000010000000010101000000001100010000;
      9'h 8e: nanoOutput = 68'b00000000000000000000000100000000010010100000001100110001011000011000;
      9'h 8f: nanoOutput = 68'b01100001000000011000000000010000100110000000011000100000001001000000;
      9'h 90: nanoOutput = 68'b00000000000000000000000000001000000100011100000001100000000001000001;
      9'h 91: nanoOutput = 68'b00010010000000000000000000010010110110000000001110000010001000011000;
      9'h 92: nanoOutput = 68'b01000001000000000000100000010010010000000000010000110001000100011000;
      9'h 93: nanoOutput = 68'b00010010000000000000010000010000110110000000001110000010001000011000;
      9'h 94: nanoOutput = 68'b01000001000000000000000010000000010100001010001000110000000001000000;
      9'h 95: nanoOutput = 68'b01000001000000000000010000001000101000000110000101000000000000110001;
      9'h 96: nanoOutput = 68'b00000001000000000000010000000000100000000000000101000100001000010000;
      9'h 97: nanoOutput = 68'b00101000000000001000010000000000000000000000000010000000000000000000;
      9'h 98: nanoOutput = 68'b00100010000000011000000000000000100000000000000010000100011000000000;
      9'h 99: nanoOutput = 68'b00100010001000011010000000000000100000000000000010000100000100000000;
      9'h 9a: nanoOutput = 68'b11010011001000000100000000010000011000010000000010000000000000000000;
      9'h 9b: nanoOutput = 68'b00010010000000000100000000000000010000000000010010001000000001000000;
      9'h 9c: nanoOutput = 68'b00001000000000011000001000000000000000000000000101110000000000000011;
      9'h 9d: nanoOutput = 68'b00100010110000000000010000001000001000000000000101000000000000110001;
      9'h 9e: nanoOutput = 68'b00100010000000011000000000000000100010100000000010000000000000000000;
      9'h 9f: nanoOutput = 68'b00100000000000011000000000110001100100011111011001100000000011000010;
      9'h a0: nanoOutput = 68'b00100000000000011000000000001000100110000000001001010000001001000001;
      9'h a1: nanoOutput = 68'b01000001000000000000000000010000000100000000011100100000000001011000;
      9'h a2: nanoOutput = 68'b00000000100000000010100000000000000001000000000101000000100000010000;
      9'h a3: nanoOutput = 68'b00000001000000000000000000011001000100000000011001000000000011000001;
      9'h a4: nanoOutput = 68'b00000000011000000010100001000110000101000000000000010000100101010000;
      9'h a5: nanoOutput = 68'b00100001000000011100000001011001000100000000011001000000000011000001;
      9'h a6: nanoOutput = 68'b01000000000000000000000000000000000101001010001101100000100001000000;
      9'h a7: nanoOutput = 68'b00000000000100000000000000000000100001001010000101100100100100010000;
      9'h a8: nanoOutput = 68'b00000000011000000000000000000010110110000000001100000000001101011000;
      9'h a9: nanoOutput = 68'b01000001000000000000000000000001111001100000001010000000110010100000;
      9'h aa: nanoOutput = 68'b00110010000000011000000000010010100010000000001110000010001000011000;
      9'h ab: nanoOutput = 68'b11000001000000000000000000011001100110110000010001000000011011000001;
      9'h ac: nanoOutput = 68'b00100000000000011010000000100001110000001100001010000000000010000010;
      9'h ad: nanoOutput = 68'b00000000000000000000000000010000000100010101010001100000000001000000;
      9'h ae: nanoOutput = 68'b01000000000000000000000000000000000010100000000010000000011000001000;
      9'h af: nanoOutput = 68'b00000001000000000000000000000000000001101010001101000000110000010000;
      9'h b0: nanoOutput = 68'b10000000000000000000001000001101100100010000000001000000000001000001;
      9'h b1: nanoOutput = 68'b01110101000000000000000000000000110000000000000010001100000101000000;
      9'h b2: nanoOutput = 68'b11000001000000000000000000001000000100010000000001000000000001000001;
      9'h b3: nanoOutput = 68'b00100010000000011000000000001001101000000010000101000010000010110001;
      9'h b4: nanoOutput = 68'b00100010000100011000000000010010100000000000000101000000000000010000;
      9'h b5: nanoOutput = 68'b11100101000000011100000000001001000100010000001001000000000011010001;
      9'h b6: nanoOutput = 68'b00100100000100111000000000000000100000000000010101100100000100010000;
      9'h b7: nanoOutput = 68'b00100010000100011000000000011010100100000000000000000000000001011001;
      9'h b8: nanoOutput = 68'b00100000000000001000001000000000100000000000000010000100000010000000;
      9'h b9: nanoOutput = 68'b00100010000000011100001000001000100100000000000001000100001001010001;
      9'h ba: nanoOutput = 68'b00010010000000000100000100000000010001000000000010000000000000000000;
      9'h bb: nanoOutput = 68'b10000000000000000000001000011101000100010000000001000000000001000001;
      9'h bc: nanoOutput = 68'b00011000000000011000001000000000100010000000000010000000000000000000;
      9'h bd: nanoOutput = 68'b01000000000000000000000000000000000100000000000001000000000001010000;
      9'h be: nanoOutput = 68'b01000000000000000000010000010000100110000000011100100000011001001000;
      9'h bf: nanoOutput = 68'b00000000001000000010001000010001010000000000000010001000000000100000;
      9'h c0: nanoOutput = 68'b11100101000000011100000000001000001000010000000101000000000000110001;
      9'h c1: nanoOutput = 68'b01000001000000000000001000010001100000000000000010000000000000000000;
      9'h c2: nanoOutput = 68'b00110100000000000000000000000000110000000000000010001100000101000000;
      9'h c3: nanoOutput = 68'b10000000000000000000001000001000100100010000010001000100000011000001;
      9'h c4: nanoOutput = 68'b01110101000000000100001000000001110000000000010010001000000001000000;
      9'h c5: nanoOutput = 68'b10000000000000000000001000001000100100010000000001000100000011000001;
      9'h c6: nanoOutput = 68'b00110100000000000000000000000000110000000000010010001100000101000000;
      9'h c7: nanoOutput = 68'b00110100000000000000000000000000110000000000010010001100011001000000;
      9'h c8: nanoOutput = 68'b01000000000000000000000000010000000110100000011100100000011001001000;
      9'h c9: nanoOutput = 68'b00000000000100000000000000010000111000000000010101000100000100110010;
      9'h ca: nanoOutput = 68'b00000000000100000000000000100010100001100000000001000000110000011000;
      9'h cb: nanoOutput = 68'b01000000000000000000000000010010000110000000010000100000001101001000;
      9'h cc: nanoOutput = 68'b00000000000000000000000000001000000110000000001001000000001001001001;
      9'h cd: nanoOutput = 68'b01000000000000000000010000000001100000000000000101000010000010010000;
      9'h ce: nanoOutput = 68'b01000000000000000000000000001000000110000000001001010000001001000001;
      9'h cf: nanoOutput = 68'b00000001000000000000000000000000000001101010001101000000110000000000;
      9'h d0: nanoOutput = 68'b11100101000000011000000000010000111001110000010010000100110100100000;
      9'h d1: nanoOutput = 68'b00000000000000000000000000011010101010000000000101000010001000110001;
      9'h d2: nanoOutput = 68'b11000001000000000000001000001101100100010000000001000000000001000001;
      9'h d3: nanoOutput = 68'b00000000000000000000000100000000010000000000000001100001000000000000;
      9'h d4: nanoOutput = 68'b00000000000000000000000000001001100100000000001001000000000011010001;
      9'h d5: nanoOutput = 68'b11000001000000000000010000010001100000010000010010000000011010000000;
      9'h d6: nanoOutput = 68'b00000000000000000000000000000000000000010110000010000000000000000000;
      9'h d7: nanoOutput = 68'b00000000000000000000000000000000000000001100000000000001000000000000;
      9'h d8: nanoOutput = 68'b00100010000000011000000000000000100010100000000010000000000000000000;
      9'h d9: nanoOutput = 68'b00001000000000011000001000000000000000000000000101110000000000000011;
      9'h da: nanoOutput = 68'b10000000000000000000000000000000000000010000000010000000000000000000;
      9'h db: nanoOutput = 68'b00000000000000000000010000000000100010000000000010000010001000000000;
      9'h dc: nanoOutput = 68'b00101000000000001000001000000000000000000000000010000000000000000000;
      9'h dd: nanoOutput = 68'b01010011000000000000100000000010100001100000001100000000110000011000;
      9'h de: nanoOutput = 68'b00000001000010000000000001000000000000000000000101000000000000010000;
      9'h df: nanoOutput = 68'b00100010000000011000010000001101101000000000000101000000000000110001;
      9'h e0: nanoOutput = 68'b00000000000000000000100000010010010000000000010000110001000100000000;
      9'h e1: nanoOutput = 68'b01000000000000000000000000010000000100000000011100100000000001000000;
      9'h e2: nanoOutput = 68'b00000000000000000000000100010010010000000000010000110001000100000000;
      9'h e3: nanoOutput = 68'b01000000000000000000100000000000010000000000000001000000110000010000;
      9'h e4: nanoOutput = 68'b01010011000000001000010000000000000001100000001100000000110000011000;
      9'h e5: nanoOutput = 68'b01000001000000000000010000001001101000000000000101000000000000110001;
      9'h e6: nanoOutput = 68'b00100100000100011001000000000000100000000000010101000100000100010000;
      9'h e7: nanoOutput = 68'b01100010000000011000100000010010110010000000001100000000110000011000;
      9'h e8: nanoOutput = 68'b00011000000000011000001000000000000000000000000101110000000000000011;
      9'h e9: nanoOutput = 68'b00000000000000000000000000001000000100000000000001000000000001010001;
      9'h ea: nanoOutput = 68'b00010010000000000100000100000000010001000000000010000000000000000000;
      9'h eb: nanoOutput = 68'b00001010000000011000001000000000000000000000000101110000000000000011;
      9'h ec: nanoOutput = 68'b00010010000000000000000000000001110100000010001110000010000010011000;
      9'h ed: nanoOutput = 68'b01100010000000011000100000010010110010000000001100000001000000011000;
      9'h ee: nanoOutput = 68'b01000000000000000000100000000010010000000000001100110001000100011000;
      9'h ef: nanoOutput = 68'b00100010000100011000000001011010100100000000000001000000000001011001;
      9'h f0: nanoOutput = 68'b00000001000000000000010000000001100001001010000101000000100000010000;
      9'h f1: nanoOutput = 68'b00000000000000000000010000000000100101000110001110000000100001011000;
      9'h f2: nanoOutput = 68'b00000000000000000000100000010010010000000000010000110001000100011000;
      9'h f3: nanoOutput = 68'b01010011000000000000100000000001100001100010001100000010110010011000;
      9'h f4: nanoOutput = 68'b01100011000000011000000000010010100100000000011101110000000001011000;
      9'h f5: nanoOutput = 68'b00000000000100000001000000010000100100000000011101000100000101010000;
      9'h f6: nanoOutput = 68'b00100010000100011000000001010010100100000000011100010000000001010000;
      9'h f7: nanoOutput = 68'b00000001000000000000010000000000100000000001000101000100000010010000;
      9'h f8: nanoOutput = 68'b00000001000000000000010000000001100000001111000101000000000000010000;
      9'h f9: nanoOutput = 68'b00000000000000000000000000010010100000000110010101100000000100000000;
      9'h fa: nanoOutput = 68'b00000111000000000000010000010000111000001000010110000100001000100000;
      9'h fb: nanoOutput = 68'b01000000000000000000100000000001110000000000001001000000110010010000;
      9'h fc: nanoOutput = 68'b01001011000000011000001000000000000001100000000000000000110000000000;
      9'h fd: nanoOutput = 68'b00000000000000000000010000000000100010000000000101000000000000010000;
      9'h fe: nanoOutput = 68'b10100100000000011100000000001000000100010000000001000000000001000001;
      9'h ff: nanoOutput = 68'b00010000000000000000000000010000100100000010000010000000000000000000;
      9'h100: nanoOutput = 68'b00000000000000000000000000001000000100000010000000110010000001000001;
      9'h101: nanoOutput = 68'b01000000000000000000000000001001100100000000001001010000000011000001;
      9'h102: nanoOutput = 68'b00000000000000000000000000001001100100000000001001010000000011000001;
      9'h103: nanoOutput = 68'b00100000000000011000000000010010100010000000010101000000001100010000;
      9'h104: nanoOutput = 68'b00000000000100000000000000000000101000000000000101000100011000110000;
      9'h105: nanoOutput = 68'b00000000000100100000100000010010010000000000010000110001000100011000;
      9'h106: nanoOutput = 68'b01000000000000000000010000010001100000000000010101000010000010010000;
      9'h107: nanoOutput = 68'b00100001000000011100010100000000110010000000001110001000100000011000;
      9'h108: nanoOutput = 68'b00000000000000000000001000000000100000000110000101000000000000000000;
      9'h109: nanoOutput = 68'b00000110000000000000000000000000000000001000000010000000000000000000;
      9'h10a: nanoOutput = 68'b01000000000000000000010000000000100100001010001100110010000001000000;
      9'h10b: nanoOutput = 68'b01000000000000000000000000000000000100001010001100000000000001000000;
      9'h10c: nanoOutput = 68'b01100001000000011000000000000000100001100010000000000000110000000000;
      9'h10d: nanoOutput = 68'b01000001000000000000010000000000100000000110000101010000000000010000;
      9'h10e: nanoOutput = 68'b00101000000000001000010000001000101010000000000101100000000000100001;
      9'h10f: nanoOutput = 68'b10000110000000000000000000001000001000001000000101100000000000100001;
      9'h110: nanoOutput = 68'b00000000000000000000000000001000000100000000000001000000000001010001;
      9'h111: nanoOutput = 68'b00100010000100111000100000000000110010100000000001000000110000010000;
      9'h112: nanoOutput = 68'b00100100000100111100000000001000000100000000000001000000000001011001;
      9'h113: nanoOutput = 68'b00100011000000011000010100000000010000000000001110001000100000011000;
      9'h114: nanoOutput = 68'b00000000000000000000000000011001100110100000010001000000011011010001;
      9'h115: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h116: nanoOutput = 68'b00000000000100100000010001001000100100000000000001000000011001001001;
      9'h117: nanoOutput = 68'b00100100001000111100001000000000100010000000000101000000000000010000;
      9'h118: nanoOutput = 68'b01000001000000000000000000010001100000000010000010000000000000000000;
      9'h119: nanoOutput = 68'b00100010000000011010000000000000110100000000011110001100100100011000;
      9'h11a: nanoOutput = 68'b11100101000000011100000100000000001000010000010101000000011010000000;
      9'h11b: nanoOutput = 68'b00010000000000000000100000000000100001100010001100000000110000000000;
      9'h11c: nanoOutput = 68'b00100010000100111000010001001000000100000000000000000000000001011001;
      9'h11d: nanoOutput = 68'b00010000000000000010000000000000100100000010001110000000000000011000;
      9'h11e: nanoOutput = 68'b11100011000000011100001000010101100000010000000101000000000000000000;
      9'h11f: nanoOutput = 68'b00100000000000011000000000110010100100011111010001100000000001000000;
      9'h120: nanoOutput = 68'b10000000000100000000000000001000100110110000000001000000000001011001;
      9'h121: nanoOutput = 68'b11000001000000000000000000001001000100010000001001000000000011010001;
      9'h122: nanoOutput = 68'b00100100000100111100000000000000000000000000000101100000000000010000;
      9'h123: nanoOutput = 68'b10000000000100100000000001001001000100010000001001000000000011001001;
      9'h124: nanoOutput = 68'b11000001000000000000000000000000000000010000000010000000000000000000;
      9'h125: nanoOutput = 68'b00110100001100100000000000000000100000000000000101100100000100010000;
      9'h126: nanoOutput = 68'b00000001000001000000000001000000000000000000000101000000000000010000;
      9'h127: nanoOutput = 68'b00000001000010000000010001000000100000000000000101000100000010010000;
      9'h128: nanoOutput = 68'b00100000000100111000000000010000101000010111010101000100000100110010;
      9'h129: nanoOutput = 68'b11100101000000011100000000000000000000010000000010000000000000000000;
      9'h12a: nanoOutput = 68'b11100101000000011000000000000000100000010000010010000100000100000000;
      9'h12b: nanoOutput = 68'b00000000000000000000000000001000001000000000000101000000000000110001;
      9'h12c: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h12d: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h12e: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h12f: nanoOutput = 68'b00000001000000000000000000001000001001100000000001000000110000110001;
      9'h130: nanoOutput = 68'b00000001000001000000000001001000000100000000000001010000000001011001;
      9'h131: nanoOutput = 68'b00100000000000001000001000000000100000000000000010000100000010000000;
      9'h132: nanoOutput = 68'b11000001000000000000010000001001001000010000000101000000000000110001;
      9'h133: nanoOutput = 68'b00000000000110000000000001000000100000000000000101000100000100010000;
      9'h134: nanoOutput = 68'b00000000000101000000000001000000100000000000000101000100000100010000;
      9'h135: nanoOutput = 68'b00000000000010100000000001010000000100000000000101000000000000010000;
      9'h136: nanoOutput = 68'b00000000000101000000000001001010000100000000000001010000000001011001;
      9'h137: nanoOutput = 68'b11100101001000011100000000000000010000010000010010001000000000100000;
      9'h138: nanoOutput = 68'b00100000000000001000000000001000001000000000000110000000000000110001;
      9'h139: nanoOutput = 68'b00100000000000011000000000000000100000000100011100000101000100011000;
      9'h13a: nanoOutput = 68'b00100000000000011000000000010000110100000000011100000101000100011000;
      9'h13b: nanoOutput = 68'b01100011100000011000000100010010000000000000000101110000000000000011;
      9'h13c: nanoOutput = 68'b01100010000000011000010100000000010000000000001100000001000000011000;
      9'h13d: nanoOutput = 68'b10000000000100100000000001001000000100010000000001000000000001011001;
      9'h13e: nanoOutput = 68'b01100010000000011000010100000010010000000000001100110001000100011000;
      9'h13f: nanoOutput = 68'b01100011000000011000010000010000000100000000011101110000000001011000;
      9'h140: nanoOutput = 68'b00000000000000000000010000000000100000000110000101000000000000010000;
      9'h141: nanoOutput = 68'b00000000000000000000000000000000000000011100001110000000000000011000;
      9'h142: nanoOutput = 68'b10100000000000001000010000001000101000000110000101000000000000100001;
      9'h143: nanoOutput = 68'b00100000000000011000000000110001100100001111011001100000000011000010;
      9'h144: nanoOutput = 68'b00000001000000000000010000000001100001001010000101000010100010010000;
      9'h145: nanoOutput = 68'b00100010001000111000010000010000000100000000011101000000000001010000;
      9'h146: nanoOutput = 68'b00100100000100111100000000000000000000000000000101000000000000010000;
      9'h147: nanoOutput = 68'b00100010000100011000010001010000000100000000011100010000000001010000;
      9'h148: nanoOutput = 68'b01000001000000000000000100010000011000000000000010000000000000000000;
      9'h149: nanoOutput = 68'b00000000000000000000010000000000100010000000000101000010001000010000;
      9'h14a: nanoOutput = 68'b00100000000100111000000000000000100000000010000100100000000000010000;
      9'h14b: nanoOutput = 68'b00100010000000011000010000001000001000000000000101000000000000110001;
      9'h14c: nanoOutput = 68'b00000001000000000000010000000000100000000000000101000100000010010000;
      9'h14d: nanoOutput = 68'b00000000000000000000000000000000000000000000000010000000000000000000;
      9'h14e: nanoOutput = 68'b00000000000000000000001000000000100100000000000000110010000001011000;
      9'h14f: nanoOutput = 68'b00000000011000000000000000000010110110000000001100000000001101011000;
    endcase
  end
endmodule
