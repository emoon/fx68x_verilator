// Produced from .sv files

module fx68k_case_box(in_0, out_0);
  input [7:0] in_0;
  output [136:0] out_0;
  wire [7:0] in_0;
  wire [136:0] out_0;
  wire n_9, n_12, n_13, n_15, n_16, n_17, n_19, n_20;
  wire n_21, n_23, n_25, n_31, n_32, n_33, n_34, n_35;
  wire n_37, n_38, n_40, n_42, n_44, n_49, n_50, n_51;
  wire n_52, n_54, n_56, n_58, n_60, n_65, n_66, n_68;
  wire n_70, n_71, n_73, n_79, n_80, n_81, n_83, n_84;
  wire n_86, n_88, n_90, n_91, n_92, n_101, n_114, n_116;
  wire n_118, n_120, n_122, n_123, n_125, n_126, n_128, n_130;
  wire n_140, n_141, n_142, n_147, n_160, n_161, n_166, n_179;
  wire n_180, n_185, n_198, n_200, n_202, n_204, n_2322, n_2323;
  wire n_2324;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[136], n_2324, n_13);
  nand g2 (n_2324, n_2322, n_2323);
  not g3 (n_2322, in_0[3]);
  nor g4 (n_2323, in_0[6], in_0[2]);
  nand g5 (n_13, n_9, n_12);
  nor g6 (n_9, in_0[1], in_0[5]);
  nor g7 (n_12, in_0[0], in_0[4]);
  nor g8 (out_0[135], n_2324, n_17);
  nand g9 (n_17, n_9, n_16);
  nor g10 (n_16, n_15, in_0[4]);
  not g11 (n_15, in_0[0]);
  nor g12 (out_0[134], n_2324, n_21);
  nand g13 (n_21, n_12, n_20);
  nor g14 (n_20, n_19, in_0[5]);
  not g15 (n_19, in_0[1]);
  nor g16 (out_0[133], n_2324, n_23);
  nand g17 (n_23, n_20, n_16);
  nor g18 (out_0[132], n_13, n_25);
  nand g19 (n_25, n_2323, in_0[3]);
  nor g20 (out_0[131], n_17, n_25);
  nor g21 (out_0[130], n_21, n_25);
  nor g22 (out_0[129], n_23, n_25);
  nor g23 (out_0[128], n_32, n_35);
  nand g24 (n_32, n_2322, n_31);
  nor g25 (n_31, in_0[7], in_0[2]);
  nand g26 (n_35, n_9, n_34);
  nor g27 (n_34, in_0[0], n_33);
  not g28 (n_33, in_0[4]);
  nor g29 (out_0[127], n_32, n_38);
  nand g30 (n_38, n_9, n_37);
  nor g31 (n_37, n_15, n_33);
  nor g32 (out_0[126], n_32, n_40);
  nand g33 (n_40, n_20, n_34);
  nor g34 (out_0[125], n_32, n_42);
  nand g35 (n_42, n_20, n_37);
  nor g36 (out_0[124], n_35, n_44);
  nand g37 (n_44, n_31, in_0[3]);
  nor g38 (out_0[123], n_38, n_44);
  nor g39 (out_0[122], n_40, n_44);
  nor g40 (out_0[121], n_42, n_44);
  nor g41 (out_0[120], n_51, n_52);
  nand g42 (n_51, n_2322, n_50);
  nor g43 (n_50, in_0[7], n_49);
  not g44 (n_49, in_0[5]);
  nand g45 (n_52, n_12, n_19);
  nor g46 (out_0[119], n_51, n_54);
  nand g47 (n_54, n_16, n_19);
  nor g48 (out_0[118], n_51, n_56);
  nand g49 (n_56, n_12, in_0[1]);
  nor g50 (out_0[117], n_51, n_58);
  nand g51 (n_58, n_16, in_0[1]);
  nor g52 (out_0[116], n_52, n_60);
  nand g53 (n_60, n_50, in_0[3]);
  nor g54 (out_0[115], n_60, n_54);
  nor g55 (out_0[114], n_60, n_56);
  nor g56 (out_0[113], n_60, n_58);
  nor g57 (out_0[112], n_2324, n_66);
  nand g58 (n_66, n_34, n_65);
  nor g59 (n_65, in_0[1], n_49);
  nor g60 (out_0[111], n_2324, n_68);
  nand g61 (n_68, n_65, n_37);
  nor g62 (out_0[110], n_2324, n_71);
  nand g63 (n_71, n_34, n_70);
  nor g64 (n_70, n_19, n_49);
  nor g65 (out_0[109], n_2324, n_73);
  nand g66 (n_73, n_70, n_37);
  nor g67 (out_0[108], n_66, n_25);
  nor g68 (out_0[107], n_68, n_25);
  nor g69 (out_0[106], n_71, n_25);
  nor g70 (out_0[105], n_73, n_25);
  nor g71 (out_0[104], n_32, n_81);
  nand g72 (n_81, n_9, n_80);
  nor g73 (n_80, in_0[0], n_79);
  not g74 (n_79, in_0[6]);
  nor g75 (out_0[103], n_32, n_84);
  nand g76 (n_84, n_9, n_83);
  nor g77 (n_83, n_15, n_79);
  nor g78 (out_0[102], n_32, n_86);
  nand g79 (n_86, n_20, n_80);
  nor g80 (out_0[101], n_32, n_88);
  nand g81 (n_88, n_20, n_83);
  nor g82 (out_0[100], n_52, n_92);
  nand g83 (n_92, n_2322, n_91);
  nor g84 (n_91, in_0[7], n_90);
  not g85 (n_90, in_0[2]);
  nor g86 (out_0[99], n_92, n_54);
  nor g87 (out_0[98], n_92, n_56);
  nor g88 (out_0[97], n_92, n_58);
  nor g89 (out_0[96], n_81, n_44);
  nor g90 (out_0[95], n_84, n_44);
  nor g91 (out_0[94], n_86, n_44);
  nor g92 (out_0[93], n_88, n_44);
  nor g93 (out_0[92], n_52, n_101);
  nand g94 (n_101, n_91, in_0[3]);
  nor g95 (out_0[91], n_101, n_54);
  nor g96 (out_0[90], n_101, n_56);
  nor g97 (out_0[89], n_101, n_58);
  nor g98 (out_0[88], n_35, n_92);
  nor g99 (out_0[87], n_38, n_92);
  nor g100 (out_0[86], n_40, n_92);
  nor g101 (out_0[85], n_42, n_92);
  nor g102 (out_0[84], n_35, n_101);
  nor g103 (out_0[83], n_38, n_101);
  nor g104 (out_0[82], n_40, n_101);
  nor g105 (out_0[81], n_42, n_101);
  nor g106 (out_0[80], n_32, n_114);
  nand g107 (n_114, n_65, n_80);
  nor g108 (out_0[79], n_32, n_116);
  nand g109 (n_116, n_65, n_83);
  nor g110 (out_0[78], n_32, n_118);
  nand g111 (n_118, n_70, n_80);
  nor g112 (out_0[77], n_32, n_120);
  nand g113 (n_120, n_70, n_83);
  nor g114 (out_0[76], n_51, n_123);
  nand g115 (n_123, n_19, n_122);
  nor g116 (n_122, in_0[0], n_90);
  nor g117 (out_0[75], n_51, n_126);
  nand g118 (n_126, n_19, n_125);
  nor g119 (n_125, n_15, n_90);
  nor g120 (out_0[74], n_51, n_128);
  nand g121 (n_128, n_122, in_0[1]);
  nor g122 (out_0[73], n_51, n_130);
  nand g123 (n_130, n_125, in_0[1]);
  nor g124 (out_0[72], n_114, n_44);
  nor g125 (out_0[71], n_116, n_44);
  nor g126 (out_0[70], n_118, n_44);
  nor g127 (out_0[69], n_120, n_44);
  nor g128 (out_0[68], n_60, n_123);
  nor g129 (out_0[67], n_60, n_126);
  nor g130 (out_0[66], n_60, n_128);
  nor g131 (out_0[65], n_60, n_130);
  nor g132 (out_0[64], n_13, n_142);
  nand g133 (n_142, n_2322, n_141);
  nor g134 (n_141, n_140, n_90);
  not g135 (n_140, in_0[7]);
  nor g136 (out_0[63], n_17, n_142);
  nor g137 (out_0[62], n_21, n_142);
  nor g138 (out_0[61], n_23, n_142);
  nor g139 (out_0[60], n_13, n_147);
  nand g140 (n_147, n_141, in_0[3]);
  nor g141 (out_0[59], n_17, n_147);
  nor g142 (out_0[58], n_21, n_147);
  nor g143 (out_0[57], n_23, n_147);
  nor g144 (out_0[56], n_35, n_142);
  nor g145 (out_0[55], n_38, n_142);
  nor g146 (out_0[54], n_40, n_142);
  nor g147 (out_0[53], n_42, n_142);
  nor g148 (out_0[52], n_35, n_147);
  nor g149 (out_0[51], n_38, n_147);
  nor g150 (out_0[50], n_40, n_147);
  nor g151 (out_0[49], n_42, n_147);
  nor g152 (out_0[48], n_123, n_161);
  nand g153 (n_161, n_2322, n_160);
  nor g154 (n_160, in_0[4], n_49);
  nor g155 (out_0[47], n_161, n_126);
  nor g156 (out_0[46], n_161, n_128);
  nor g157 (out_0[45], n_161, n_130);
  nor g158 (out_0[44], n_123, n_166);
  nand g159 (n_166, n_160, in_0[3]);
  nor g160 (out_0[43], n_166, n_126);
  nor g161 (out_0[42], n_166, n_128);
  nor g162 (out_0[41], n_166, n_130);
  nor g163 (out_0[40], n_66, n_142);
  nor g164 (out_0[39], n_68, n_142);
  nor g165 (out_0[38], n_71, n_142);
  nor g166 (out_0[37], n_73, n_142);
  nor g167 (out_0[36], n_66, n_147);
  nor g168 (out_0[35], n_68, n_147);
  nor g169 (out_0[34], n_71, n_147);
  nor g170 (out_0[33], n_73, n_147);
  nor g171 (out_0[32], n_13, n_180);
  nand g172 (n_180, n_2322, n_179);
  nor g173 (n_179, n_140, in_0[2]);
  nor g174 (out_0[31], n_17, n_180);
  nor g175 (out_0[30], n_21, n_180);
  nor g176 (out_0[29], n_23, n_180);
  nor g177 (out_0[28], n_13, n_185);
  nand g178 (n_185, n_179, in_0[3]);
  nor g179 (out_0[27], n_17, n_185);
  nor g180 (out_0[26], n_21, n_185);
  nor g181 (out_0[25], n_23, n_185);
  nor g182 (out_0[24], n_35, n_180);
  nor g183 (out_0[23], n_38, n_180);
  nor g184 (out_0[22], n_40, n_180);
  nor g185 (out_0[21], n_42, n_180);
  nor g186 (out_0[20], n_35, n_185);
  nor g187 (out_0[19], n_38, n_185);
  nor g188 (out_0[18], n_40, n_185);
  nor g189 (out_0[17], n_42, n_185);
  nor g190 (out_0[16], n_180, n_198);
  nand g191 (n_198, n_65, n_12);
  nor g192 (out_0[15], n_180, n_200);
  nand g193 (n_200, n_65, n_16);
  nor g194 (out_0[14], n_180, n_202);
  nand g195 (n_202, n_70, n_12);
  nor g196 (out_0[13], n_180, n_204);
  nand g197 (n_204, n_70, n_16);
  nor g198 (out_0[12], n_198, n_185);
  nor g199 (out_0[11], n_200, n_185);
  nor g200 (out_0[10], n_202, n_185);
  nor g201 (out_0[9], n_204, n_185);
  nor g202 (out_0[8], n_66, n_180);
  nor g203 (out_0[7], n_68, n_180);
  nor g204 (out_0[6], n_71, n_180);
  nor g205 (out_0[5], n_73, n_180);
  nor g206 (out_0[4], n_66, n_185);
  nor g207 (out_0[3], n_68, n_185);
  nor g208 (out_0[2], n_71, n_185);
  nor g209 (out_0[1], n_73, n_185);
endmodule

module fx68k_mux(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7,
     in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16,
     in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25,
     in_26, in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34,
     in_35, in_36, in_37, in_38, in_39, in_40, in_41, in_42, in_43,
     in_44, in_45, in_46, in_47, in_48, in_49, in_50, in_51, in_52,
     in_53, in_54, in_55, in_56, in_57, in_58, in_59, in_60, in_61,
     in_62, in_63, in_64, in_65, in_66, in_67, in_68, in_69, in_70,
     in_71, in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79,
     in_80, in_81, in_82, in_83, in_84, in_85, in_86, in_87, in_88,
     in_89, in_90, in_91, in_92, in_93, in_94, in_95, in_96, in_97,
     in_98, in_99, in_100, in_101, in_102, in_103, in_104, in_105,
     in_106, in_107, in_108, in_109, in_110, in_111, in_112, in_113,
     in_114, in_115, in_116, in_117, in_118, in_119, in_120, in_121,
     in_122, in_123, in_124, in_125, in_126, in_127, in_128, in_129,
     in_130, in_131, in_132, in_133, in_134, in_135, z);
  input [135:0] ctl;
  input [6:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17,
       in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26,
       in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35,
       in_36, in_37, in_38, in_39, in_40, in_41, in_42, in_43, in_44,
       in_45, in_46, in_47, in_48, in_49, in_50, in_51, in_52, in_53,
       in_54, in_55, in_56, in_57, in_58, in_59, in_60, in_61, in_62,
       in_63, in_64, in_65, in_66, in_67, in_68, in_69, in_70, in_71,
       in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, in_80,
       in_81, in_82, in_83, in_84, in_85, in_86, in_87, in_88, in_89,
       in_90, in_91, in_92, in_93, in_94, in_95, in_96, in_97, in_98,
       in_99, in_100, in_101, in_102, in_103, in_104, in_105, in_106,
       in_107, in_108, in_109, in_110, in_111, in_112, in_113, in_114,
       in_115, in_116, in_117, in_118, in_119, in_120, in_121, in_122,
       in_123, in_124, in_125, in_126, in_127, in_128, in_129, in_130,
       in_131, in_132, in_133, in_134, in_135;
  output [6:0] z;
  wire [135:0] ctl;
  wire [6:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17,
       in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26,
       in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35,
       in_36, in_37, in_38, in_39, in_40, in_41, in_42, in_43, in_44,
       in_45, in_46, in_47, in_48, in_49, in_50, in_51, in_52, in_53,
       in_54, in_55, in_56, in_57, in_58, in_59, in_60, in_61, in_62,
       in_63, in_64, in_65, in_66, in_67, in_68, in_69, in_70, in_71,
       in_72, in_73, in_74, in_75, in_76, in_77, in_78, in_79, in_80,
       in_81, in_82, in_83, in_84, in_85, in_86, in_87, in_88, in_89,
       in_90, in_91, in_92, in_93, in_94, in_95, in_96, in_97, in_98,
       in_99, in_100, in_101, in_102, in_103, in_104, in_105, in_106,
       in_107, in_108, in_109, in_110, in_111, in_112, in_113, in_114,
       in_115, in_116, in_117, in_118, in_119, in_120, in_121, in_122,
       in_123, in_124, in_125, in_126, in_127, in_128, in_129, in_130,
       in_131, in_132, in_133, in_134, in_135;
  wire [6:0] z;
  CDN_mux136 g1(.sel0 (ctl[135]), .data0 (in_0[6]), .sel1 (ctl[134]),
       .data1 (in_1[6]), .sel2 (ctl[133]), .data2 (in_2[6]), .sel3
       (ctl[132]), .data3 (in_3[6]), .sel4 (ctl[131]), .data4
       (in_4[6]), .sel5 (ctl[130]), .data5 (in_5[6]), .sel6 (ctl[129]),
       .data6 (in_6[6]), .sel7 (ctl[128]), .data7 (in_7[6]), .sel8
       (ctl[127]), .data8 (in_8[6]), .sel9 (ctl[126]), .data9
       (in_9[6]), .sel10 (ctl[125]), .data10 (in_10[6]), .sel11
       (ctl[124]), .data11 (in_11[6]), .sel12 (ctl[123]), .data12
       (in_12[6]), .sel13 (ctl[122]), .data13 (in_13[6]), .sel14
       (ctl[121]), .data14 (in_14[6]), .sel15 (ctl[120]), .data15
       (in_15[6]), .sel16 (ctl[119]), .data16 (in_16[6]), .sel17
       (ctl[118]), .data17 (in_17[6]), .sel18 (ctl[117]), .data18
       (in_18[6]), .sel19 (ctl[116]), .data19 (in_19[6]), .sel20
       (ctl[115]), .data20 (in_20[6]), .sel21 (ctl[114]), .data21
       (in_21[6]), .sel22 (ctl[113]), .data22 (in_22[6]), .sel23
       (ctl[112]), .data23 (in_23[6]), .sel24 (ctl[111]), .data24
       (in_24[6]), .sel25 (ctl[110]), .data25 (in_25[6]), .sel26
       (ctl[109]), .data26 (in_26[6]), .sel27 (ctl[108]), .data27
       (in_27[6]), .sel28 (ctl[107]), .data28 (in_28[6]), .sel29
       (ctl[106]), .data29 (in_29[6]), .sel30 (ctl[105]), .data30
       (in_30[6]), .sel31 (ctl[104]), .data31 (in_31[6]), .sel32
       (ctl[103]), .data32 (in_32[6]), .sel33 (ctl[102]), .data33
       (in_33[6]), .sel34 (ctl[101]), .data34 (in_34[6]), .sel35
       (ctl[100]), .data35 (in_35[6]), .sel36 (ctl[99]), .data36
       (in_36[6]), .sel37 (ctl[98]), .data37 (in_37[6]), .sel38
       (ctl[97]), .data38 (in_38[6]), .sel39 (ctl[96]), .data39
       (in_39[6]), .sel40 (ctl[95]), .data40 (in_40[6]), .sel41
       (ctl[94]), .data41 (in_41[6]), .sel42 (ctl[93]), .data42
       (in_42[6]), .sel43 (ctl[92]), .data43 (in_43[6]), .sel44
       (ctl[91]), .data44 (in_44[6]), .sel45 (ctl[90]), .data45
       (in_45[6]), .sel46 (ctl[89]), .data46 (in_46[6]), .sel47
       (ctl[88]), .data47 (in_47[6]), .sel48 (ctl[87]), .data48
       (in_48[6]), .sel49 (ctl[86]), .data49 (in_49[6]), .sel50
       (ctl[85]), .data50 (in_50[6]), .sel51 (ctl[84]), .data51
       (in_51[6]), .sel52 (ctl[83]), .data52 (in_52[6]), .sel53
       (ctl[82]), .data53 (in_53[6]), .sel54 (ctl[81]), .data54
       (in_54[6]), .sel55 (ctl[80]), .data55 (in_55[6]), .sel56
       (ctl[79]), .data56 (in_56[6]), .sel57 (ctl[78]), .data57
       (in_57[6]), .sel58 (ctl[77]), .data58 (in_58[6]), .sel59
       (ctl[76]), .data59 (in_59[6]), .sel60 (ctl[75]), .data60
       (in_60[6]), .sel61 (ctl[74]), .data61 (in_61[6]), .sel62
       (ctl[73]), .data62 (in_62[6]), .sel63 (ctl[72]), .data63
       (in_63[6]), .sel64 (ctl[71]), .data64 (in_64[6]), .sel65
       (ctl[70]), .data65 (in_65[6]), .sel66 (ctl[69]), .data66
       (in_66[6]), .sel67 (ctl[68]), .data67 (in_67[6]), .sel68
       (ctl[67]), .data68 (in_68[6]), .sel69 (ctl[66]), .data69
       (in_69[6]), .sel70 (ctl[65]), .data70 (in_70[6]), .sel71
       (ctl[64]), .data71 (in_71[6]), .sel72 (ctl[63]), .data72
       (in_72[6]), .sel73 (ctl[62]), .data73 (in_73[6]), .sel74
       (ctl[61]), .data74 (in_74[6]), .sel75 (ctl[60]), .data75
       (in_75[6]), .sel76 (ctl[59]), .data76 (in_76[6]), .sel77
       (ctl[58]), .data77 (in_77[6]), .sel78 (ctl[57]), .data78
       (in_78[6]), .sel79 (ctl[56]), .data79 (in_79[6]), .sel80
       (ctl[55]), .data80 (in_80[6]), .sel81 (ctl[54]), .data81
       (in_81[6]), .sel82 (ctl[53]), .data82 (in_82[6]), .sel83
       (ctl[52]), .data83 (in_83[6]), .sel84 (ctl[51]), .data84
       (in_84[6]), .sel85 (ctl[50]), .data85 (in_85[6]), .sel86
       (ctl[49]), .data86 (in_86[6]), .sel87 (ctl[48]), .data87
       (in_87[6]), .sel88 (ctl[47]), .data88 (in_88[6]), .sel89
       (ctl[46]), .data89 (in_89[6]), .sel90 (ctl[45]), .data90
       (in_90[6]), .sel91 (ctl[44]), .data91 (in_91[6]), .sel92
       (ctl[43]), .data92 (in_92[6]), .sel93 (ctl[42]), .data93
       (in_93[6]), .sel94 (ctl[41]), .data94 (in_94[6]), .sel95
       (ctl[40]), .data95 (in_95[6]), .sel96 (ctl[39]), .data96
       (in_96[6]), .sel97 (ctl[38]), .data97 (in_97[6]), .sel98
       (ctl[37]), .data98 (in_98[6]), .sel99 (ctl[36]), .data99
       (in_99[6]), .sel100 (ctl[35]), .data100 (in_100[6]), .sel101
       (ctl[34]), .data101 (in_101[6]), .sel102 (ctl[33]), .data102
       (in_102[6]), .sel103 (ctl[32]), .data103 (in_103[6]), .sel104
       (ctl[31]), .data104 (in_104[6]), .sel105 (ctl[30]), .data105
       (in_105[6]), .sel106 (ctl[29]), .data106 (in_106[6]), .sel107
       (ctl[28]), .data107 (in_107[6]), .sel108 (ctl[27]), .data108
       (in_108[6]), .sel109 (ctl[26]), .data109 (in_109[6]), .sel110
       (ctl[25]), .data110 (in_110[6]), .sel111 (ctl[24]), .data111
       (in_111[6]), .sel112 (ctl[23]), .data112 (in_112[6]), .sel113
       (ctl[22]), .data113 (in_113[6]), .sel114 (ctl[21]), .data114
       (in_114[6]), .sel115 (ctl[20]), .data115 (in_115[6]), .sel116
       (ctl[19]), .data116 (in_116[6]), .sel117 (ctl[18]), .data117
       (in_117[6]), .sel118 (ctl[17]), .data118 (in_118[6]), .sel119
       (ctl[16]), .data119 (in_119[6]), .sel120 (ctl[15]), .data120
       (in_120[6]), .sel121 (ctl[14]), .data121 (in_121[6]), .sel122
       (ctl[13]), .data122 (in_122[6]), .sel123 (ctl[12]), .data123
       (in_123[6]), .sel124 (ctl[11]), .data124 (in_124[6]), .sel125
       (ctl[10]), .data125 (in_125[6]), .sel126 (ctl[9]), .data126
       (in_126[6]), .sel127 (ctl[8]), .data127 (in_127[6]), .sel128
       (ctl[7]), .data128 (in_128[6]), .sel129 (ctl[6]), .data129
       (in_129[6]), .sel130 (ctl[5]), .data130 (in_130[6]), .sel131
       (ctl[4]), .data131 (in_131[6]), .sel132 (ctl[3]), .data132
       (in_132[6]), .sel133 (ctl[2]), .data133 (in_133[6]), .sel134
       (ctl[1]), .data134 (in_134[6]), .sel135 (ctl[0]), .data135
       (in_135[6]), .z (z[6]));
  CDN_mux136 g8(.sel0 (ctl[135]), .data0 (in_0[5]), .sel1 (ctl[134]),
       .data1 (in_1[5]), .sel2 (ctl[133]), .data2 (in_2[5]), .sel3
       (ctl[132]), .data3 (in_3[5]), .sel4 (ctl[131]), .data4
       (in_4[5]), .sel5 (ctl[130]), .data5 (in_5[5]), .sel6 (ctl[129]),
       .data6 (in_6[5]), .sel7 (ctl[128]), .data7 (in_7[5]), .sel8
       (ctl[127]), .data8 (in_8[5]), .sel9 (ctl[126]), .data9
       (in_9[5]), .sel10 (ctl[125]), .data10 (in_10[5]), .sel11
       (ctl[124]), .data11 (in_11[5]), .sel12 (ctl[123]), .data12
       (in_12[5]), .sel13 (ctl[122]), .data13 (in_13[5]), .sel14
       (ctl[121]), .data14 (in_14[5]), .sel15 (ctl[120]), .data15
       (in_15[5]), .sel16 (ctl[119]), .data16 (in_16[5]), .sel17
       (ctl[118]), .data17 (in_17[5]), .sel18 (ctl[117]), .data18
       (in_18[5]), .sel19 (ctl[116]), .data19 (in_19[5]), .sel20
       (ctl[115]), .data20 (in_20[5]), .sel21 (ctl[114]), .data21
       (in_21[5]), .sel22 (ctl[113]), .data22 (in_22[5]), .sel23
       (ctl[112]), .data23 (in_23[5]), .sel24 (ctl[111]), .data24
       (in_24[5]), .sel25 (ctl[110]), .data25 (in_25[5]), .sel26
       (ctl[109]), .data26 (in_26[5]), .sel27 (ctl[108]), .data27
       (in_27[5]), .sel28 (ctl[107]), .data28 (in_28[5]), .sel29
       (ctl[106]), .data29 (in_29[5]), .sel30 (ctl[105]), .data30
       (in_30[5]), .sel31 (ctl[104]), .data31 (in_31[5]), .sel32
       (ctl[103]), .data32 (in_32[5]), .sel33 (ctl[102]), .data33
       (in_33[5]), .sel34 (ctl[101]), .data34 (in_34[5]), .sel35
       (ctl[100]), .data35 (in_35[5]), .sel36 (ctl[99]), .data36
       (in_36[5]), .sel37 (ctl[98]), .data37 (in_37[5]), .sel38
       (ctl[97]), .data38 (in_38[5]), .sel39 (ctl[96]), .data39
       (in_39[5]), .sel40 (ctl[95]), .data40 (in_40[5]), .sel41
       (ctl[94]), .data41 (in_41[5]), .sel42 (ctl[93]), .data42
       (in_42[5]), .sel43 (ctl[92]), .data43 (in_43[5]), .sel44
       (ctl[91]), .data44 (in_44[5]), .sel45 (ctl[90]), .data45
       (in_45[5]), .sel46 (ctl[89]), .data46 (in_46[5]), .sel47
       (ctl[88]), .data47 (in_47[5]), .sel48 (ctl[87]), .data48
       (in_48[5]), .sel49 (ctl[86]), .data49 (in_49[5]), .sel50
       (ctl[85]), .data50 (in_50[5]), .sel51 (ctl[84]), .data51
       (in_51[5]), .sel52 (ctl[83]), .data52 (in_52[5]), .sel53
       (ctl[82]), .data53 (in_53[5]), .sel54 (ctl[81]), .data54
       (in_54[5]), .sel55 (ctl[80]), .data55 (in_55[5]), .sel56
       (ctl[79]), .data56 (in_56[5]), .sel57 (ctl[78]), .data57
       (in_57[5]), .sel58 (ctl[77]), .data58 (in_58[5]), .sel59
       (ctl[76]), .data59 (in_59[5]), .sel60 (ctl[75]), .data60
       (in_60[5]), .sel61 (ctl[74]), .data61 (in_61[5]), .sel62
       (ctl[73]), .data62 (in_62[5]), .sel63 (ctl[72]), .data63
       (in_63[5]), .sel64 (ctl[71]), .data64 (in_64[5]), .sel65
       (ctl[70]), .data65 (in_65[5]), .sel66 (ctl[69]), .data66
       (in_66[5]), .sel67 (ctl[68]), .data67 (in_67[5]), .sel68
       (ctl[67]), .data68 (in_68[5]), .sel69 (ctl[66]), .data69
       (in_69[5]), .sel70 (ctl[65]), .data70 (in_70[5]), .sel71
       (ctl[64]), .data71 (in_71[5]), .sel72 (ctl[63]), .data72
       (in_72[5]), .sel73 (ctl[62]), .data73 (in_73[5]), .sel74
       (ctl[61]), .data74 (in_74[5]), .sel75 (ctl[60]), .data75
       (in_75[5]), .sel76 (ctl[59]), .data76 (in_76[5]), .sel77
       (ctl[58]), .data77 (in_77[5]), .sel78 (ctl[57]), .data78
       (in_78[5]), .sel79 (ctl[56]), .data79 (in_79[5]), .sel80
       (ctl[55]), .data80 (in_80[5]), .sel81 (ctl[54]), .data81
       (in_81[5]), .sel82 (ctl[53]), .data82 (in_82[5]), .sel83
       (ctl[52]), .data83 (in_83[5]), .sel84 (ctl[51]), .data84
       (in_84[5]), .sel85 (ctl[50]), .data85 (in_85[5]), .sel86
       (ctl[49]), .data86 (in_86[5]), .sel87 (ctl[48]), .data87
       (in_87[5]), .sel88 (ctl[47]), .data88 (in_88[5]), .sel89
       (ctl[46]), .data89 (in_89[5]), .sel90 (ctl[45]), .data90
       (in_90[5]), .sel91 (ctl[44]), .data91 (in_91[5]), .sel92
       (ctl[43]), .data92 (in_92[5]), .sel93 (ctl[42]), .data93
       (in_93[5]), .sel94 (ctl[41]), .data94 (in_94[5]), .sel95
       (ctl[40]), .data95 (in_95[5]), .sel96 (ctl[39]), .data96
       (in_96[5]), .sel97 (ctl[38]), .data97 (in_97[5]), .sel98
       (ctl[37]), .data98 (in_98[5]), .sel99 (ctl[36]), .data99
       (in_99[5]), .sel100 (ctl[35]), .data100 (in_100[5]), .sel101
       (ctl[34]), .data101 (in_101[5]), .sel102 (ctl[33]), .data102
       (in_102[5]), .sel103 (ctl[32]), .data103 (in_103[5]), .sel104
       (ctl[31]), .data104 (in_104[5]), .sel105 (ctl[30]), .data105
       (in_105[5]), .sel106 (ctl[29]), .data106 (in_106[5]), .sel107
       (ctl[28]), .data107 (in_107[5]), .sel108 (ctl[27]), .data108
       (in_108[5]), .sel109 (ctl[26]), .data109 (in_109[5]), .sel110
       (ctl[25]), .data110 (in_110[5]), .sel111 (ctl[24]), .data111
       (in_111[5]), .sel112 (ctl[23]), .data112 (in_112[5]), .sel113
       (ctl[22]), .data113 (in_113[5]), .sel114 (ctl[21]), .data114
       (in_114[5]), .sel115 (ctl[20]), .data115 (in_115[5]), .sel116
       (ctl[19]), .data116 (in_116[5]), .sel117 (ctl[18]), .data117
       (in_117[5]), .sel118 (ctl[17]), .data118 (in_118[5]), .sel119
       (ctl[16]), .data119 (in_119[5]), .sel120 (ctl[15]), .data120
       (in_120[5]), .sel121 (ctl[14]), .data121 (in_121[5]), .sel122
       (ctl[13]), .data122 (in_122[5]), .sel123 (ctl[12]), .data123
       (in_123[5]), .sel124 (ctl[11]), .data124 (in_124[5]), .sel125
       (ctl[10]), .data125 (in_125[5]), .sel126 (ctl[9]), .data126
       (in_126[5]), .sel127 (ctl[8]), .data127 (in_127[5]), .sel128
       (ctl[7]), .data128 (in_128[5]), .sel129 (ctl[6]), .data129
       (in_129[5]), .sel130 (ctl[5]), .data130 (in_130[5]), .sel131
       (ctl[4]), .data131 (in_131[5]), .sel132 (ctl[3]), .data132
       (in_132[5]), .sel133 (ctl[2]), .data133 (in_133[5]), .sel134
       (ctl[1]), .data134 (in_134[5]), .sel135 (ctl[0]), .data135
       (in_135[5]), .z (z[5]));
  CDN_mux136 g9(.sel0 (ctl[135]), .data0 (in_0[4]), .sel1 (ctl[134]),
       .data1 (in_1[4]), .sel2 (ctl[133]), .data2 (in_2[4]), .sel3
       (ctl[132]), .data3 (in_3[4]), .sel4 (ctl[131]), .data4
       (in_4[4]), .sel5 (ctl[130]), .data5 (in_5[4]), .sel6 (ctl[129]),
       .data6 (in_6[4]), .sel7 (ctl[128]), .data7 (in_7[4]), .sel8
       (ctl[127]), .data8 (in_8[4]), .sel9 (ctl[126]), .data9
       (in_9[4]), .sel10 (ctl[125]), .data10 (in_10[4]), .sel11
       (ctl[124]), .data11 (in_11[4]), .sel12 (ctl[123]), .data12
       (in_12[4]), .sel13 (ctl[122]), .data13 (in_13[4]), .sel14
       (ctl[121]), .data14 (in_14[4]), .sel15 (ctl[120]), .data15
       (in_15[4]), .sel16 (ctl[119]), .data16 (in_16[4]), .sel17
       (ctl[118]), .data17 (in_17[4]), .sel18 (ctl[117]), .data18
       (in_18[4]), .sel19 (ctl[116]), .data19 (in_19[4]), .sel20
       (ctl[115]), .data20 (in_20[4]), .sel21 (ctl[114]), .data21
       (in_21[4]), .sel22 (ctl[113]), .data22 (in_22[4]), .sel23
       (ctl[112]), .data23 (in_23[4]), .sel24 (ctl[111]), .data24
       (in_24[4]), .sel25 (ctl[110]), .data25 (in_25[4]), .sel26
       (ctl[109]), .data26 (in_26[4]), .sel27 (ctl[108]), .data27
       (in_27[4]), .sel28 (ctl[107]), .data28 (in_28[4]), .sel29
       (ctl[106]), .data29 (in_29[4]), .sel30 (ctl[105]), .data30
       (in_30[4]), .sel31 (ctl[104]), .data31 (in_31[4]), .sel32
       (ctl[103]), .data32 (in_32[4]), .sel33 (ctl[102]), .data33
       (in_33[4]), .sel34 (ctl[101]), .data34 (in_34[4]), .sel35
       (ctl[100]), .data35 (in_35[4]), .sel36 (ctl[99]), .data36
       (in_36[4]), .sel37 (ctl[98]), .data37 (in_37[4]), .sel38
       (ctl[97]), .data38 (in_38[4]), .sel39 (ctl[96]), .data39
       (in_39[4]), .sel40 (ctl[95]), .data40 (in_40[4]), .sel41
       (ctl[94]), .data41 (in_41[4]), .sel42 (ctl[93]), .data42
       (in_42[4]), .sel43 (ctl[92]), .data43 (in_43[4]), .sel44
       (ctl[91]), .data44 (in_44[4]), .sel45 (ctl[90]), .data45
       (in_45[4]), .sel46 (ctl[89]), .data46 (in_46[4]), .sel47
       (ctl[88]), .data47 (in_47[4]), .sel48 (ctl[87]), .data48
       (in_48[4]), .sel49 (ctl[86]), .data49 (in_49[4]), .sel50
       (ctl[85]), .data50 (in_50[4]), .sel51 (ctl[84]), .data51
       (in_51[4]), .sel52 (ctl[83]), .data52 (in_52[4]), .sel53
       (ctl[82]), .data53 (in_53[4]), .sel54 (ctl[81]), .data54
       (in_54[4]), .sel55 (ctl[80]), .data55 (in_55[4]), .sel56
       (ctl[79]), .data56 (in_56[4]), .sel57 (ctl[78]), .data57
       (in_57[4]), .sel58 (ctl[77]), .data58 (in_58[4]), .sel59
       (ctl[76]), .data59 (in_59[4]), .sel60 (ctl[75]), .data60
       (in_60[4]), .sel61 (ctl[74]), .data61 (in_61[4]), .sel62
       (ctl[73]), .data62 (in_62[4]), .sel63 (ctl[72]), .data63
       (in_63[4]), .sel64 (ctl[71]), .data64 (in_64[4]), .sel65
       (ctl[70]), .data65 (in_65[4]), .sel66 (ctl[69]), .data66
       (in_66[4]), .sel67 (ctl[68]), .data67 (in_67[4]), .sel68
       (ctl[67]), .data68 (in_68[4]), .sel69 (ctl[66]), .data69
       (in_69[4]), .sel70 (ctl[65]), .data70 (in_70[4]), .sel71
       (ctl[64]), .data71 (in_71[4]), .sel72 (ctl[63]), .data72
       (in_72[4]), .sel73 (ctl[62]), .data73 (in_73[4]), .sel74
       (ctl[61]), .data74 (in_74[4]), .sel75 (ctl[60]), .data75
       (in_75[4]), .sel76 (ctl[59]), .data76 (in_76[4]), .sel77
       (ctl[58]), .data77 (in_77[4]), .sel78 (ctl[57]), .data78
       (in_78[4]), .sel79 (ctl[56]), .data79 (in_79[4]), .sel80
       (ctl[55]), .data80 (in_80[4]), .sel81 (ctl[54]), .data81
       (in_81[4]), .sel82 (ctl[53]), .data82 (in_82[4]), .sel83
       (ctl[52]), .data83 (in_83[4]), .sel84 (ctl[51]), .data84
       (in_84[4]), .sel85 (ctl[50]), .data85 (in_85[4]), .sel86
       (ctl[49]), .data86 (in_86[4]), .sel87 (ctl[48]), .data87
       (in_87[4]), .sel88 (ctl[47]), .data88 (in_88[4]), .sel89
       (ctl[46]), .data89 (in_89[4]), .sel90 (ctl[45]), .data90
       (in_90[4]), .sel91 (ctl[44]), .data91 (in_91[4]), .sel92
       (ctl[43]), .data92 (in_92[4]), .sel93 (ctl[42]), .data93
       (in_93[4]), .sel94 (ctl[41]), .data94 (in_94[4]), .sel95
       (ctl[40]), .data95 (in_95[4]), .sel96 (ctl[39]), .data96
       (in_96[4]), .sel97 (ctl[38]), .data97 (in_97[4]), .sel98
       (ctl[37]), .data98 (in_98[4]), .sel99 (ctl[36]), .data99
       (in_99[4]), .sel100 (ctl[35]), .data100 (in_100[4]), .sel101
       (ctl[34]), .data101 (in_101[4]), .sel102 (ctl[33]), .data102
       (in_102[4]), .sel103 (ctl[32]), .data103 (in_103[4]), .sel104
       (ctl[31]), .data104 (in_104[4]), .sel105 (ctl[30]), .data105
       (in_105[4]), .sel106 (ctl[29]), .data106 (in_106[4]), .sel107
       (ctl[28]), .data107 (in_107[4]), .sel108 (ctl[27]), .data108
       (in_108[4]), .sel109 (ctl[26]), .data109 (in_109[4]), .sel110
       (ctl[25]), .data110 (in_110[4]), .sel111 (ctl[24]), .data111
       (in_111[4]), .sel112 (ctl[23]), .data112 (in_112[4]), .sel113
       (ctl[22]), .data113 (in_113[4]), .sel114 (ctl[21]), .data114
       (in_114[4]), .sel115 (ctl[20]), .data115 (in_115[4]), .sel116
       (ctl[19]), .data116 (in_116[4]), .sel117 (ctl[18]), .data117
       (in_117[4]), .sel118 (ctl[17]), .data118 (in_118[4]), .sel119
       (ctl[16]), .data119 (in_119[4]), .sel120 (ctl[15]), .data120
       (in_120[4]), .sel121 (ctl[14]), .data121 (in_121[4]), .sel122
       (ctl[13]), .data122 (in_122[4]), .sel123 (ctl[12]), .data123
       (in_123[4]), .sel124 (ctl[11]), .data124 (in_124[4]), .sel125
       (ctl[10]), .data125 (in_125[4]), .sel126 (ctl[9]), .data126
       (in_126[4]), .sel127 (ctl[8]), .data127 (in_127[4]), .sel128
       (ctl[7]), .data128 (in_128[4]), .sel129 (ctl[6]), .data129
       (in_129[4]), .sel130 (ctl[5]), .data130 (in_130[4]), .sel131
       (ctl[4]), .data131 (in_131[4]), .sel132 (ctl[3]), .data132
       (in_132[4]), .sel133 (ctl[2]), .data133 (in_133[4]), .sel134
       (ctl[1]), .data134 (in_134[4]), .sel135 (ctl[0]), .data135
       (in_135[4]), .z (z[4]));
  CDN_mux136 g10(.sel0 (ctl[135]), .data0 (in_0[3]), .sel1 (ctl[134]),
       .data1 (in_1[3]), .sel2 (ctl[133]), .data2 (in_2[3]), .sel3
       (ctl[132]), .data3 (in_3[3]), .sel4 (ctl[131]), .data4
       (in_4[3]), .sel5 (ctl[130]), .data5 (in_5[3]), .sel6 (ctl[129]),
       .data6 (in_6[3]), .sel7 (ctl[128]), .data7 (in_7[3]), .sel8
       (ctl[127]), .data8 (in_8[3]), .sel9 (ctl[126]), .data9
       (in_9[3]), .sel10 (ctl[125]), .data10 (in_10[3]), .sel11
       (ctl[124]), .data11 (in_11[3]), .sel12 (ctl[123]), .data12
       (in_12[3]), .sel13 (ctl[122]), .data13 (in_13[3]), .sel14
       (ctl[121]), .data14 (in_14[3]), .sel15 (ctl[120]), .data15
       (in_15[3]), .sel16 (ctl[119]), .data16 (in_16[3]), .sel17
       (ctl[118]), .data17 (in_17[3]), .sel18 (ctl[117]), .data18
       (in_18[3]), .sel19 (ctl[116]), .data19 (in_19[3]), .sel20
       (ctl[115]), .data20 (in_20[3]), .sel21 (ctl[114]), .data21
       (in_21[3]), .sel22 (ctl[113]), .data22 (in_22[3]), .sel23
       (ctl[112]), .data23 (in_23[3]), .sel24 (ctl[111]), .data24
       (in_24[3]), .sel25 (ctl[110]), .data25 (in_25[3]), .sel26
       (ctl[109]), .data26 (in_26[3]), .sel27 (ctl[108]), .data27
       (in_27[3]), .sel28 (ctl[107]), .data28 (in_28[3]), .sel29
       (ctl[106]), .data29 (in_29[3]), .sel30 (ctl[105]), .data30
       (in_30[3]), .sel31 (ctl[104]), .data31 (in_31[3]), .sel32
       (ctl[103]), .data32 (in_32[3]), .sel33 (ctl[102]), .data33
       (in_33[3]), .sel34 (ctl[101]), .data34 (in_34[3]), .sel35
       (ctl[100]), .data35 (in_35[3]), .sel36 (ctl[99]), .data36
       (in_36[3]), .sel37 (ctl[98]), .data37 (in_37[3]), .sel38
       (ctl[97]), .data38 (in_38[3]), .sel39 (ctl[96]), .data39
       (in_39[3]), .sel40 (ctl[95]), .data40 (in_40[3]), .sel41
       (ctl[94]), .data41 (in_41[3]), .sel42 (ctl[93]), .data42
       (in_42[3]), .sel43 (ctl[92]), .data43 (in_43[3]), .sel44
       (ctl[91]), .data44 (in_44[3]), .sel45 (ctl[90]), .data45
       (in_45[3]), .sel46 (ctl[89]), .data46 (in_46[3]), .sel47
       (ctl[88]), .data47 (in_47[3]), .sel48 (ctl[87]), .data48
       (in_48[3]), .sel49 (ctl[86]), .data49 (in_49[3]), .sel50
       (ctl[85]), .data50 (in_50[3]), .sel51 (ctl[84]), .data51
       (in_51[3]), .sel52 (ctl[83]), .data52 (in_52[3]), .sel53
       (ctl[82]), .data53 (in_53[3]), .sel54 (ctl[81]), .data54
       (in_54[3]), .sel55 (ctl[80]), .data55 (in_55[3]), .sel56
       (ctl[79]), .data56 (in_56[3]), .sel57 (ctl[78]), .data57
       (in_57[3]), .sel58 (ctl[77]), .data58 (in_58[3]), .sel59
       (ctl[76]), .data59 (in_59[3]), .sel60 (ctl[75]), .data60
       (in_60[3]), .sel61 (ctl[74]), .data61 (in_61[3]), .sel62
       (ctl[73]), .data62 (in_62[3]), .sel63 (ctl[72]), .data63
       (in_63[3]), .sel64 (ctl[71]), .data64 (in_64[3]), .sel65
       (ctl[70]), .data65 (in_65[3]), .sel66 (ctl[69]), .data66
       (in_66[3]), .sel67 (ctl[68]), .data67 (in_67[3]), .sel68
       (ctl[67]), .data68 (in_68[3]), .sel69 (ctl[66]), .data69
       (in_69[3]), .sel70 (ctl[65]), .data70 (in_70[3]), .sel71
       (ctl[64]), .data71 (in_71[3]), .sel72 (ctl[63]), .data72
       (in_72[3]), .sel73 (ctl[62]), .data73 (in_73[3]), .sel74
       (ctl[61]), .data74 (in_74[3]), .sel75 (ctl[60]), .data75
       (in_75[3]), .sel76 (ctl[59]), .data76 (in_76[3]), .sel77
       (ctl[58]), .data77 (in_77[3]), .sel78 (ctl[57]), .data78
       (in_78[3]), .sel79 (ctl[56]), .data79 (in_79[3]), .sel80
       (ctl[55]), .data80 (in_80[3]), .sel81 (ctl[54]), .data81
       (in_81[3]), .sel82 (ctl[53]), .data82 (in_82[3]), .sel83
       (ctl[52]), .data83 (in_83[3]), .sel84 (ctl[51]), .data84
       (in_84[3]), .sel85 (ctl[50]), .data85 (in_85[3]), .sel86
       (ctl[49]), .data86 (in_86[3]), .sel87 (ctl[48]), .data87
       (in_87[3]), .sel88 (ctl[47]), .data88 (in_88[3]), .sel89
       (ctl[46]), .data89 (in_89[3]), .sel90 (ctl[45]), .data90
       (in_90[3]), .sel91 (ctl[44]), .data91 (in_91[3]), .sel92
       (ctl[43]), .data92 (in_92[3]), .sel93 (ctl[42]), .data93
       (in_93[3]), .sel94 (ctl[41]), .data94 (in_94[3]), .sel95
       (ctl[40]), .data95 (in_95[3]), .sel96 (ctl[39]), .data96
       (in_96[3]), .sel97 (ctl[38]), .data97 (in_97[3]), .sel98
       (ctl[37]), .data98 (in_98[3]), .sel99 (ctl[36]), .data99
       (in_99[3]), .sel100 (ctl[35]), .data100 (in_100[3]), .sel101
       (ctl[34]), .data101 (in_101[3]), .sel102 (ctl[33]), .data102
       (in_102[3]), .sel103 (ctl[32]), .data103 (in_103[3]), .sel104
       (ctl[31]), .data104 (in_104[3]), .sel105 (ctl[30]), .data105
       (in_105[3]), .sel106 (ctl[29]), .data106 (in_106[3]), .sel107
       (ctl[28]), .data107 (in_107[3]), .sel108 (ctl[27]), .data108
       (in_108[3]), .sel109 (ctl[26]), .data109 (in_109[3]), .sel110
       (ctl[25]), .data110 (in_110[3]), .sel111 (ctl[24]), .data111
       (in_111[3]), .sel112 (ctl[23]), .data112 (in_112[3]), .sel113
       (ctl[22]), .data113 (in_113[3]), .sel114 (ctl[21]), .data114
       (in_114[3]), .sel115 (ctl[20]), .data115 (in_115[3]), .sel116
       (ctl[19]), .data116 (in_116[3]), .sel117 (ctl[18]), .data117
       (in_117[3]), .sel118 (ctl[17]), .data118 (in_118[3]), .sel119
       (ctl[16]), .data119 (in_119[3]), .sel120 (ctl[15]), .data120
       (in_120[3]), .sel121 (ctl[14]), .data121 (in_121[3]), .sel122
       (ctl[13]), .data122 (in_122[3]), .sel123 (ctl[12]), .data123
       (in_123[3]), .sel124 (ctl[11]), .data124 (in_124[3]), .sel125
       (ctl[10]), .data125 (in_125[3]), .sel126 (ctl[9]), .data126
       (in_126[3]), .sel127 (ctl[8]), .data127 (in_127[3]), .sel128
       (ctl[7]), .data128 (in_128[3]), .sel129 (ctl[6]), .data129
       (in_129[3]), .sel130 (ctl[5]), .data130 (in_130[3]), .sel131
       (ctl[4]), .data131 (in_131[3]), .sel132 (ctl[3]), .data132
       (in_132[3]), .sel133 (ctl[2]), .data133 (in_133[3]), .sel134
       (ctl[1]), .data134 (in_134[3]), .sel135 (ctl[0]), .data135
       (in_135[3]), .z (z[3]));
  CDN_mux136 g11(.sel0 (ctl[135]), .data0 (in_0[2]), .sel1 (ctl[134]),
       .data1 (in_1[2]), .sel2 (ctl[133]), .data2 (in_2[2]), .sel3
       (ctl[132]), .data3 (in_3[2]), .sel4 (ctl[131]), .data4
       (in_4[2]), .sel5 (ctl[130]), .data5 (in_5[2]), .sel6 (ctl[129]),
       .data6 (in_6[2]), .sel7 (ctl[128]), .data7 (in_7[2]), .sel8
       (ctl[127]), .data8 (in_8[2]), .sel9 (ctl[126]), .data9
       (in_9[2]), .sel10 (ctl[125]), .data10 (in_10[2]), .sel11
       (ctl[124]), .data11 (in_11[2]), .sel12 (ctl[123]), .data12
       (in_12[2]), .sel13 (ctl[122]), .data13 (in_13[2]), .sel14
       (ctl[121]), .data14 (in_14[2]), .sel15 (ctl[120]), .data15
       (in_15[2]), .sel16 (ctl[119]), .data16 (in_16[2]), .sel17
       (ctl[118]), .data17 (in_17[2]), .sel18 (ctl[117]), .data18
       (in_18[2]), .sel19 (ctl[116]), .data19 (in_19[2]), .sel20
       (ctl[115]), .data20 (in_20[2]), .sel21 (ctl[114]), .data21
       (in_21[2]), .sel22 (ctl[113]), .data22 (in_22[2]), .sel23
       (ctl[112]), .data23 (in_23[2]), .sel24 (ctl[111]), .data24
       (in_24[2]), .sel25 (ctl[110]), .data25 (in_25[2]), .sel26
       (ctl[109]), .data26 (in_26[2]), .sel27 (ctl[108]), .data27
       (in_27[2]), .sel28 (ctl[107]), .data28 (in_28[2]), .sel29
       (ctl[106]), .data29 (in_29[2]), .sel30 (ctl[105]), .data30
       (in_30[2]), .sel31 (ctl[104]), .data31 (in_31[2]), .sel32
       (ctl[103]), .data32 (in_32[2]), .sel33 (ctl[102]), .data33
       (in_33[2]), .sel34 (ctl[101]), .data34 (in_34[2]), .sel35
       (ctl[100]), .data35 (in_35[2]), .sel36 (ctl[99]), .data36
       (in_36[2]), .sel37 (ctl[98]), .data37 (in_37[2]), .sel38
       (ctl[97]), .data38 (in_38[2]), .sel39 (ctl[96]), .data39
       (in_39[2]), .sel40 (ctl[95]), .data40 (in_40[2]), .sel41
       (ctl[94]), .data41 (in_41[2]), .sel42 (ctl[93]), .data42
       (in_42[2]), .sel43 (ctl[92]), .data43 (in_43[2]), .sel44
       (ctl[91]), .data44 (in_44[2]), .sel45 (ctl[90]), .data45
       (in_45[2]), .sel46 (ctl[89]), .data46 (in_46[2]), .sel47
       (ctl[88]), .data47 (in_47[2]), .sel48 (ctl[87]), .data48
       (in_48[2]), .sel49 (ctl[86]), .data49 (in_49[2]), .sel50
       (ctl[85]), .data50 (in_50[2]), .sel51 (ctl[84]), .data51
       (in_51[2]), .sel52 (ctl[83]), .data52 (in_52[2]), .sel53
       (ctl[82]), .data53 (in_53[2]), .sel54 (ctl[81]), .data54
       (in_54[2]), .sel55 (ctl[80]), .data55 (in_55[2]), .sel56
       (ctl[79]), .data56 (in_56[2]), .sel57 (ctl[78]), .data57
       (in_57[2]), .sel58 (ctl[77]), .data58 (in_58[2]), .sel59
       (ctl[76]), .data59 (in_59[2]), .sel60 (ctl[75]), .data60
       (in_60[2]), .sel61 (ctl[74]), .data61 (in_61[2]), .sel62
       (ctl[73]), .data62 (in_62[2]), .sel63 (ctl[72]), .data63
       (in_63[2]), .sel64 (ctl[71]), .data64 (in_64[2]), .sel65
       (ctl[70]), .data65 (in_65[2]), .sel66 (ctl[69]), .data66
       (in_66[2]), .sel67 (ctl[68]), .data67 (in_67[2]), .sel68
       (ctl[67]), .data68 (in_68[2]), .sel69 (ctl[66]), .data69
       (in_69[2]), .sel70 (ctl[65]), .data70 (in_70[2]), .sel71
       (ctl[64]), .data71 (in_71[2]), .sel72 (ctl[63]), .data72
       (in_72[2]), .sel73 (ctl[62]), .data73 (in_73[2]), .sel74
       (ctl[61]), .data74 (in_74[2]), .sel75 (ctl[60]), .data75
       (in_75[2]), .sel76 (ctl[59]), .data76 (in_76[2]), .sel77
       (ctl[58]), .data77 (in_77[2]), .sel78 (ctl[57]), .data78
       (in_78[2]), .sel79 (ctl[56]), .data79 (in_79[2]), .sel80
       (ctl[55]), .data80 (in_80[2]), .sel81 (ctl[54]), .data81
       (in_81[2]), .sel82 (ctl[53]), .data82 (in_82[2]), .sel83
       (ctl[52]), .data83 (in_83[2]), .sel84 (ctl[51]), .data84
       (in_84[2]), .sel85 (ctl[50]), .data85 (in_85[2]), .sel86
       (ctl[49]), .data86 (in_86[2]), .sel87 (ctl[48]), .data87
       (in_87[2]), .sel88 (ctl[47]), .data88 (in_88[2]), .sel89
       (ctl[46]), .data89 (in_89[2]), .sel90 (ctl[45]), .data90
       (in_90[2]), .sel91 (ctl[44]), .data91 (in_91[2]), .sel92
       (ctl[43]), .data92 (in_92[2]), .sel93 (ctl[42]), .data93
       (in_93[2]), .sel94 (ctl[41]), .data94 (in_94[2]), .sel95
       (ctl[40]), .data95 (in_95[2]), .sel96 (ctl[39]), .data96
       (in_96[2]), .sel97 (ctl[38]), .data97 (in_97[2]), .sel98
       (ctl[37]), .data98 (in_98[2]), .sel99 (ctl[36]), .data99
       (in_99[2]), .sel100 (ctl[35]), .data100 (in_100[2]), .sel101
       (ctl[34]), .data101 (in_101[2]), .sel102 (ctl[33]), .data102
       (in_102[2]), .sel103 (ctl[32]), .data103 (in_103[2]), .sel104
       (ctl[31]), .data104 (in_104[2]), .sel105 (ctl[30]), .data105
       (in_105[2]), .sel106 (ctl[29]), .data106 (in_106[2]), .sel107
       (ctl[28]), .data107 (in_107[2]), .sel108 (ctl[27]), .data108
       (in_108[2]), .sel109 (ctl[26]), .data109 (in_109[2]), .sel110
       (ctl[25]), .data110 (in_110[2]), .sel111 (ctl[24]), .data111
       (in_111[2]), .sel112 (ctl[23]), .data112 (in_112[2]), .sel113
       (ctl[22]), .data113 (in_113[2]), .sel114 (ctl[21]), .data114
       (in_114[2]), .sel115 (ctl[20]), .data115 (in_115[2]), .sel116
       (ctl[19]), .data116 (in_116[2]), .sel117 (ctl[18]), .data117
       (in_117[2]), .sel118 (ctl[17]), .data118 (in_118[2]), .sel119
       (ctl[16]), .data119 (in_119[2]), .sel120 (ctl[15]), .data120
       (in_120[2]), .sel121 (ctl[14]), .data121 (in_121[2]), .sel122
       (ctl[13]), .data122 (in_122[2]), .sel123 (ctl[12]), .data123
       (in_123[2]), .sel124 (ctl[11]), .data124 (in_124[2]), .sel125
       (ctl[10]), .data125 (in_125[2]), .sel126 (ctl[9]), .data126
       (in_126[2]), .sel127 (ctl[8]), .data127 (in_127[2]), .sel128
       (ctl[7]), .data128 (in_128[2]), .sel129 (ctl[6]), .data129
       (in_129[2]), .sel130 (ctl[5]), .data130 (in_130[2]), .sel131
       (ctl[4]), .data131 (in_131[2]), .sel132 (ctl[3]), .data132
       (in_132[2]), .sel133 (ctl[2]), .data133 (in_133[2]), .sel134
       (ctl[1]), .data134 (in_134[2]), .sel135 (ctl[0]), .data135
       (in_135[2]), .z (z[2]));
  CDN_mux136 g12(.sel0 (ctl[135]), .data0 (in_0[1]), .sel1 (ctl[134]),
       .data1 (in_1[1]), .sel2 (ctl[133]), .data2 (in_2[1]), .sel3
       (ctl[132]), .data3 (in_3[1]), .sel4 (ctl[131]), .data4
       (in_4[1]), .sel5 (ctl[130]), .data5 (in_5[1]), .sel6 (ctl[129]),
       .data6 (in_6[1]), .sel7 (ctl[128]), .data7 (in_7[1]), .sel8
       (ctl[127]), .data8 (in_8[1]), .sel9 (ctl[126]), .data9
       (in_9[1]), .sel10 (ctl[125]), .data10 (in_10[1]), .sel11
       (ctl[124]), .data11 (in_11[1]), .sel12 (ctl[123]), .data12
       (in_12[1]), .sel13 (ctl[122]), .data13 (in_13[1]), .sel14
       (ctl[121]), .data14 (in_14[1]), .sel15 (ctl[120]), .data15
       (in_15[1]), .sel16 (ctl[119]), .data16 (in_16[1]), .sel17
       (ctl[118]), .data17 (in_17[1]), .sel18 (ctl[117]), .data18
       (in_18[1]), .sel19 (ctl[116]), .data19 (in_19[1]), .sel20
       (ctl[115]), .data20 (in_20[1]), .sel21 (ctl[114]), .data21
       (in_21[1]), .sel22 (ctl[113]), .data22 (in_22[1]), .sel23
       (ctl[112]), .data23 (in_23[1]), .sel24 (ctl[111]), .data24
       (in_24[1]), .sel25 (ctl[110]), .data25 (in_25[1]), .sel26
       (ctl[109]), .data26 (in_26[1]), .sel27 (ctl[108]), .data27
       (in_27[1]), .sel28 (ctl[107]), .data28 (in_28[1]), .sel29
       (ctl[106]), .data29 (in_29[1]), .sel30 (ctl[105]), .data30
       (in_30[1]), .sel31 (ctl[104]), .data31 (in_31[1]), .sel32
       (ctl[103]), .data32 (in_32[1]), .sel33 (ctl[102]), .data33
       (in_33[1]), .sel34 (ctl[101]), .data34 (in_34[1]), .sel35
       (ctl[100]), .data35 (in_35[1]), .sel36 (ctl[99]), .data36
       (in_36[1]), .sel37 (ctl[98]), .data37 (in_37[1]), .sel38
       (ctl[97]), .data38 (in_38[1]), .sel39 (ctl[96]), .data39
       (in_39[1]), .sel40 (ctl[95]), .data40 (in_40[1]), .sel41
       (ctl[94]), .data41 (in_41[1]), .sel42 (ctl[93]), .data42
       (in_42[1]), .sel43 (ctl[92]), .data43 (in_43[1]), .sel44
       (ctl[91]), .data44 (in_44[1]), .sel45 (ctl[90]), .data45
       (in_45[1]), .sel46 (ctl[89]), .data46 (in_46[1]), .sel47
       (ctl[88]), .data47 (in_47[1]), .sel48 (ctl[87]), .data48
       (in_48[1]), .sel49 (ctl[86]), .data49 (in_49[1]), .sel50
       (ctl[85]), .data50 (in_50[1]), .sel51 (ctl[84]), .data51
       (in_51[1]), .sel52 (ctl[83]), .data52 (in_52[1]), .sel53
       (ctl[82]), .data53 (in_53[1]), .sel54 (ctl[81]), .data54
       (in_54[1]), .sel55 (ctl[80]), .data55 (in_55[1]), .sel56
       (ctl[79]), .data56 (in_56[1]), .sel57 (ctl[78]), .data57
       (in_57[1]), .sel58 (ctl[77]), .data58 (in_58[1]), .sel59
       (ctl[76]), .data59 (in_59[1]), .sel60 (ctl[75]), .data60
       (in_60[1]), .sel61 (ctl[74]), .data61 (in_61[1]), .sel62
       (ctl[73]), .data62 (in_62[1]), .sel63 (ctl[72]), .data63
       (in_63[1]), .sel64 (ctl[71]), .data64 (in_64[1]), .sel65
       (ctl[70]), .data65 (in_65[1]), .sel66 (ctl[69]), .data66
       (in_66[1]), .sel67 (ctl[68]), .data67 (in_67[1]), .sel68
       (ctl[67]), .data68 (in_68[1]), .sel69 (ctl[66]), .data69
       (in_69[1]), .sel70 (ctl[65]), .data70 (in_70[1]), .sel71
       (ctl[64]), .data71 (in_71[1]), .sel72 (ctl[63]), .data72
       (in_72[1]), .sel73 (ctl[62]), .data73 (in_73[1]), .sel74
       (ctl[61]), .data74 (in_74[1]), .sel75 (ctl[60]), .data75
       (in_75[1]), .sel76 (ctl[59]), .data76 (in_76[1]), .sel77
       (ctl[58]), .data77 (in_77[1]), .sel78 (ctl[57]), .data78
       (in_78[1]), .sel79 (ctl[56]), .data79 (in_79[1]), .sel80
       (ctl[55]), .data80 (in_80[1]), .sel81 (ctl[54]), .data81
       (in_81[1]), .sel82 (ctl[53]), .data82 (in_82[1]), .sel83
       (ctl[52]), .data83 (in_83[1]), .sel84 (ctl[51]), .data84
       (in_84[1]), .sel85 (ctl[50]), .data85 (in_85[1]), .sel86
       (ctl[49]), .data86 (in_86[1]), .sel87 (ctl[48]), .data87
       (in_87[1]), .sel88 (ctl[47]), .data88 (in_88[1]), .sel89
       (ctl[46]), .data89 (in_89[1]), .sel90 (ctl[45]), .data90
       (in_90[1]), .sel91 (ctl[44]), .data91 (in_91[1]), .sel92
       (ctl[43]), .data92 (in_92[1]), .sel93 (ctl[42]), .data93
       (in_93[1]), .sel94 (ctl[41]), .data94 (in_94[1]), .sel95
       (ctl[40]), .data95 (in_95[1]), .sel96 (ctl[39]), .data96
       (in_96[1]), .sel97 (ctl[38]), .data97 (in_97[1]), .sel98
       (ctl[37]), .data98 (in_98[1]), .sel99 (ctl[36]), .data99
       (in_99[1]), .sel100 (ctl[35]), .data100 (in_100[1]), .sel101
       (ctl[34]), .data101 (in_101[1]), .sel102 (ctl[33]), .data102
       (in_102[1]), .sel103 (ctl[32]), .data103 (in_103[1]), .sel104
       (ctl[31]), .data104 (in_104[1]), .sel105 (ctl[30]), .data105
       (in_105[1]), .sel106 (ctl[29]), .data106 (in_106[1]), .sel107
       (ctl[28]), .data107 (in_107[1]), .sel108 (ctl[27]), .data108
       (in_108[1]), .sel109 (ctl[26]), .data109 (in_109[1]), .sel110
       (ctl[25]), .data110 (in_110[1]), .sel111 (ctl[24]), .data111
       (in_111[1]), .sel112 (ctl[23]), .data112 (in_112[1]), .sel113
       (ctl[22]), .data113 (in_113[1]), .sel114 (ctl[21]), .data114
       (in_114[1]), .sel115 (ctl[20]), .data115 (in_115[1]), .sel116
       (ctl[19]), .data116 (in_116[1]), .sel117 (ctl[18]), .data117
       (in_117[1]), .sel118 (ctl[17]), .data118 (in_118[1]), .sel119
       (ctl[16]), .data119 (in_119[1]), .sel120 (ctl[15]), .data120
       (in_120[1]), .sel121 (ctl[14]), .data121 (in_121[1]), .sel122
       (ctl[13]), .data122 (in_122[1]), .sel123 (ctl[12]), .data123
       (in_123[1]), .sel124 (ctl[11]), .data124 (in_124[1]), .sel125
       (ctl[10]), .data125 (in_125[1]), .sel126 (ctl[9]), .data126
       (in_126[1]), .sel127 (ctl[8]), .data127 (in_127[1]), .sel128
       (ctl[7]), .data128 (in_128[1]), .sel129 (ctl[6]), .data129
       (in_129[1]), .sel130 (ctl[5]), .data130 (in_130[1]), .sel131
       (ctl[4]), .data131 (in_131[1]), .sel132 (ctl[3]), .data132
       (in_132[1]), .sel133 (ctl[2]), .data133 (in_133[1]), .sel134
       (ctl[1]), .data134 (in_134[1]), .sel135 (ctl[0]), .data135
       (in_135[1]), .z (z[1]));
  CDN_mux136 g13(.sel0 (ctl[135]), .data0 (in_0[0]), .sel1 (ctl[134]),
       .data1 (in_1[0]), .sel2 (ctl[133]), .data2 (in_2[0]), .sel3
       (ctl[132]), .data3 (in_3[0]), .sel4 (ctl[131]), .data4
       (in_4[0]), .sel5 (ctl[130]), .data5 (in_5[0]), .sel6 (ctl[129]),
       .data6 (in_6[0]), .sel7 (ctl[128]), .data7 (in_7[0]), .sel8
       (ctl[127]), .data8 (in_8[0]), .sel9 (ctl[126]), .data9
       (in_9[0]), .sel10 (ctl[125]), .data10 (in_10[0]), .sel11
       (ctl[124]), .data11 (in_11[0]), .sel12 (ctl[123]), .data12
       (in_12[0]), .sel13 (ctl[122]), .data13 (in_13[0]), .sel14
       (ctl[121]), .data14 (in_14[0]), .sel15 (ctl[120]), .data15
       (in_15[0]), .sel16 (ctl[119]), .data16 (in_16[0]), .sel17
       (ctl[118]), .data17 (in_17[0]), .sel18 (ctl[117]), .data18
       (in_18[0]), .sel19 (ctl[116]), .data19 (in_19[0]), .sel20
       (ctl[115]), .data20 (in_20[0]), .sel21 (ctl[114]), .data21
       (in_21[0]), .sel22 (ctl[113]), .data22 (in_22[0]), .sel23
       (ctl[112]), .data23 (in_23[0]), .sel24 (ctl[111]), .data24
       (in_24[0]), .sel25 (ctl[110]), .data25 (in_25[0]), .sel26
       (ctl[109]), .data26 (in_26[0]), .sel27 (ctl[108]), .data27
       (in_27[0]), .sel28 (ctl[107]), .data28 (in_28[0]), .sel29
       (ctl[106]), .data29 (in_29[0]), .sel30 (ctl[105]), .data30
       (in_30[0]), .sel31 (ctl[104]), .data31 (in_31[0]), .sel32
       (ctl[103]), .data32 (in_32[0]), .sel33 (ctl[102]), .data33
       (in_33[0]), .sel34 (ctl[101]), .data34 (in_34[0]), .sel35
       (ctl[100]), .data35 (in_35[0]), .sel36 (ctl[99]), .data36
       (in_36[0]), .sel37 (ctl[98]), .data37 (in_37[0]), .sel38
       (ctl[97]), .data38 (in_38[0]), .sel39 (ctl[96]), .data39
       (in_39[0]), .sel40 (ctl[95]), .data40 (in_40[0]), .sel41
       (ctl[94]), .data41 (in_41[0]), .sel42 (ctl[93]), .data42
       (in_42[0]), .sel43 (ctl[92]), .data43 (in_43[0]), .sel44
       (ctl[91]), .data44 (in_44[0]), .sel45 (ctl[90]), .data45
       (in_45[0]), .sel46 (ctl[89]), .data46 (in_46[0]), .sel47
       (ctl[88]), .data47 (in_47[0]), .sel48 (ctl[87]), .data48
       (in_48[0]), .sel49 (ctl[86]), .data49 (in_49[0]), .sel50
       (ctl[85]), .data50 (in_50[0]), .sel51 (ctl[84]), .data51
       (in_51[0]), .sel52 (ctl[83]), .data52 (in_52[0]), .sel53
       (ctl[82]), .data53 (in_53[0]), .sel54 (ctl[81]), .data54
       (in_54[0]), .sel55 (ctl[80]), .data55 (in_55[0]), .sel56
       (ctl[79]), .data56 (in_56[0]), .sel57 (ctl[78]), .data57
       (in_57[0]), .sel58 (ctl[77]), .data58 (in_58[0]), .sel59
       (ctl[76]), .data59 (in_59[0]), .sel60 (ctl[75]), .data60
       (in_60[0]), .sel61 (ctl[74]), .data61 (in_61[0]), .sel62
       (ctl[73]), .data62 (in_62[0]), .sel63 (ctl[72]), .data63
       (in_63[0]), .sel64 (ctl[71]), .data64 (in_64[0]), .sel65
       (ctl[70]), .data65 (in_65[0]), .sel66 (ctl[69]), .data66
       (in_66[0]), .sel67 (ctl[68]), .data67 (in_67[0]), .sel68
       (ctl[67]), .data68 (in_68[0]), .sel69 (ctl[66]), .data69
       (in_69[0]), .sel70 (ctl[65]), .data70 (in_70[0]), .sel71
       (ctl[64]), .data71 (in_71[0]), .sel72 (ctl[63]), .data72
       (in_72[0]), .sel73 (ctl[62]), .data73 (in_73[0]), .sel74
       (ctl[61]), .data74 (in_74[0]), .sel75 (ctl[60]), .data75
       (in_75[0]), .sel76 (ctl[59]), .data76 (in_76[0]), .sel77
       (ctl[58]), .data77 (in_77[0]), .sel78 (ctl[57]), .data78
       (in_78[0]), .sel79 (ctl[56]), .data79 (in_79[0]), .sel80
       (ctl[55]), .data80 (in_80[0]), .sel81 (ctl[54]), .data81
       (in_81[0]), .sel82 (ctl[53]), .data82 (in_82[0]), .sel83
       (ctl[52]), .data83 (in_83[0]), .sel84 (ctl[51]), .data84
       (in_84[0]), .sel85 (ctl[50]), .data85 (in_85[0]), .sel86
       (ctl[49]), .data86 (in_86[0]), .sel87 (ctl[48]), .data87
       (in_87[0]), .sel88 (ctl[47]), .data88 (in_88[0]), .sel89
       (ctl[46]), .data89 (in_89[0]), .sel90 (ctl[45]), .data90
       (in_90[0]), .sel91 (ctl[44]), .data91 (in_91[0]), .sel92
       (ctl[43]), .data92 (in_92[0]), .sel93 (ctl[42]), .data93
       (in_93[0]), .sel94 (ctl[41]), .data94 (in_94[0]), .sel95
       (ctl[40]), .data95 (in_95[0]), .sel96 (ctl[39]), .data96
       (in_96[0]), .sel97 (ctl[38]), .data97 (in_97[0]), .sel98
       (ctl[37]), .data98 (in_98[0]), .sel99 (ctl[36]), .data99
       (in_99[0]), .sel100 (ctl[35]), .data100 (in_100[0]), .sel101
       (ctl[34]), .data101 (in_101[0]), .sel102 (ctl[33]), .data102
       (in_102[0]), .sel103 (ctl[32]), .data103 (in_103[0]), .sel104
       (ctl[31]), .data104 (in_104[0]), .sel105 (ctl[30]), .data105
       (in_105[0]), .sel106 (ctl[29]), .data106 (in_106[0]), .sel107
       (ctl[28]), .data107 (in_107[0]), .sel108 (ctl[27]), .data108
       (in_108[0]), .sel109 (ctl[26]), .data109 (in_109[0]), .sel110
       (ctl[25]), .data110 (in_110[0]), .sel111 (ctl[24]), .data111
       (in_111[0]), .sel112 (ctl[23]), .data112 (in_112[0]), .sel113
       (ctl[22]), .data113 (in_113[0]), .sel114 (ctl[21]), .data114
       (in_114[0]), .sel115 (ctl[20]), .data115 (in_115[0]), .sel116
       (ctl[19]), .data116 (in_116[0]), .sel117 (ctl[18]), .data117
       (in_117[0]), .sel118 (ctl[17]), .data118 (in_118[0]), .sel119
       (ctl[16]), .data119 (in_119[0]), .sel120 (ctl[15]), .data120
       (in_120[0]), .sel121 (ctl[14]), .data121 (in_121[0]), .sel122
       (ctl[13]), .data122 (in_122[0]), .sel123 (ctl[12]), .data123
       (in_123[0]), .sel124 (ctl[11]), .data124 (in_124[0]), .sel125
       (ctl[10]), .data125 (in_125[0]), .sel126 (ctl[9]), .data126
       (in_126[0]), .sel127 (ctl[8]), .data127 (in_127[0]), .sel128
       (ctl[7]), .data128 (in_128[0]), .sel129 (ctl[6]), .data129
       (in_129[0]), .sel130 (ctl[5]), .data130 (in_130[0]), .sel131
       (ctl[4]), .data131 (in_131[0]), .sel132 (ctl[3]), .data132
       (in_132[0]), .sel133 (ctl[2]), .data133 (in_133[0]), .sel134
       (ctl[1]), .data134 (in_134[0]), .sel135 (ctl[0]), .data135
       (in_135[0]), .z (z[0]));
endmodule

module fx68k_microToNanoAddr(uAddr, orgAddr);
  input [9:0] uAddr;
  output [8:0] orgAddr;
  wire [9:0] uAddr;
  wire [8:0] orgAddr;
  wire UNCONNECTED, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967;
  wire n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975;
  wire n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983;
  wire n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991;
  wire n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999;
  wire n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007;
  wire n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031;
  wire n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039;
  wire n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047;
  wire n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055;
  wire n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063;
  wire n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071;
  wire n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079;
  wire n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087;
  wire n_1088;
  assign orgAddr[0] = uAddr[0];
  assign orgAddr[1] = uAddr[1];
  fx68k_case_box ctl_baseAddr_2479_9(.in_0 (uAddr[9:2]), .out_0
       ({n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961,
       n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970,
       n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979,
       n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988,
       n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997,
       n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005,
       n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013,
       n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021,
       n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029,
       n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037,
       n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045,
       n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053,
       n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061,
       n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069,
       n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077,
       n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085,
       n_1086, n_1087, n_1088, UNCONNECTED}));
  fx68k_mux mux_orgBase_2479_9(.ctl ({n_953, n_954, n_955, n_956,
       n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965,
       n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974,
       n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983,
       n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992,
       n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001,
       n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009,
       n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017,
       n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025,
       n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033,
       n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041,
       n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049,
       n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057,
       n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065,
       n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073,
       n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081,
       n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088}), .in_0
       (7'b0000000), .in_1 (7'b0000001), .in_2 (7'b0000010), .in_3
       (7'b0000010), .in_4 (7'b0000011), .in_5 (7'b0000100), .in_6
       (7'b0000101), .in_7 (7'b0000101), .in_8 (7'b0000110), .in_9
       (7'b0000111), .in_10 (7'b0001000), .in_11 (7'b0001000), .in_12
       (7'b0001001), .in_13 (7'b0001010), .in_14 (7'b0001011), .in_15
       (7'b0001011), .in_16 (7'b0001100), .in_17 (7'b0001101), .in_18
       (7'b0001110), .in_19 (7'b0001101), .in_20 (7'b0001111), .in_21
       (7'b0010000), .in_22 (7'b0010001), .in_23 (7'b0010000), .in_24
       (7'b0010010), .in_25 (7'b0010011), .in_26 (7'b0010100), .in_27
       (7'b0010100), .in_28 (7'b0010101), .in_29 (7'b0010110), .in_30
       (7'b0010111), .in_31 (7'b0010111), .in_32 (7'b0011000), .in_33
       (7'b0011000), .in_34 (7'b0011000), .in_35 (7'b0011000), .in_36
       (7'b0011001), .in_37 (7'b0011001), .in_38 (7'b0011001), .in_39
       (7'b0011001), .in_40 (7'b0011010), .in_41 (7'b0011010), .in_42
       (7'b0011010), .in_43 (7'b0011010), .in_44 (7'b0011011), .in_45
       (7'b0011011), .in_46 (7'b0011011), .in_47 (7'b0011011), .in_48
       (7'b0011100), .in_49 (7'b0011101), .in_50 (7'b0011110), .in_51
       (7'b0011111), .in_52 (7'b0100000), .in_53 (7'b0100001), .in_54
       (7'b0100010), .in_55 (7'b0100011), .in_56 (7'b0100100), .in_57
       (7'b0100100), .in_58 (7'b0100100), .in_59 (7'b0100100), .in_60
       (7'b0100100), .in_61 (7'b0100100), .in_62 (7'b0100100), .in_63
       (7'b0100100), .in_64 (7'b0100101), .in_65 (7'b0100101), .in_66
       (7'b0100101), .in_67 (7'b0100101), .in_68 (7'b0100101), .in_69
       (7'b0100101), .in_70 (7'b0100101), .in_71 (7'b0100101), .in_72
       (7'b0100110), .in_73 (7'b0100111), .in_74 (7'b0101000), .in_75
       (7'b0101001), .in_76 (7'b0101010), .in_77 (7'b0101011), .in_78
       (7'b0101100), .in_79 (7'b0101101), .in_80 (7'b0101110), .in_81
       (7'b0101111), .in_82 (7'b0110000), .in_83 (7'b0110001), .in_84
       (7'b0110010), .in_85 (7'b0110011), .in_86 (7'b0110100), .in_87
       (7'b0110101), .in_88 (7'b0110110), .in_89 (7'b0110110), .in_90
       (7'b0110111), .in_91 (7'b0110111), .in_92 (7'b0111000), .in_93
       (7'b0111000), .in_94 (7'b0111001), .in_95 (7'b0111001), .in_96
       (7'b0111010), .in_97 (7'b0111010), .in_98 (7'b0111011), .in_99
       (7'b0111011), .in_100 (7'b0111100), .in_101 (7'b0111100),
       .in_102 (7'b0111101), .in_103 (7'b0111101), .in_104
       (7'b0111110), .in_105 (7'b0111111), .in_106 (7'b1000000),
       .in_107 (7'b1000001), .in_108 (7'b1000010), .in_109
       (7'b1000011), .in_110 (7'b1000100), .in_111 (7'b1000101),
       .in_112 (7'b1000110), .in_113 (7'b1000111), .in_114
       (7'b1001000), .in_115 (7'b1001001), .in_116 (7'b1001010),
       .in_117 (7'b1001011), .in_118 (7'b1001100), .in_119
       (7'b1001101), .in_120 (7'b1001110), .in_121 (7'b1001110),
       .in_122 (7'b1001111), .in_123 (7'b1001111), .in_124
       (7'b1010000), .in_125 (7'b1010000), .in_126 (7'b1010001),
       .in_127 (7'b1010001), .in_128 (7'b1010010), .in_129
       (7'b1010010), .in_130 (7'b1010010), .in_131 (7'b1010010),
       .in_132 (7'b1010011), .in_133 (7'b1010011), .in_134
       (7'b1010011), .in_135 (7'b1010011), .z (orgAddr[8:2]));
endmodule

module fx68k_onehotEncoder4(bin, bitMap);
  input [3:0] bin;
  output [15:0] bitMap;
  wire [3:0] bin;
  wire [15:0] bitMap;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380;
  nand g1 (n_365, n_361, n_362, n_363, n_364);
  nand g2 (n_366, n_361, n_362, n_363, bin[0]);
  nand g3 (n_367, n_361, n_362, bin[1], n_364);
  nand g4 (n_368, n_361, n_362, bin[1], bin[0]);
  nand g5 (n_369, n_361, bin[2], n_363, n_364);
  nand g6 (n_370, n_361, bin[2], n_363, bin[0]);
  nand g7 (n_371, n_361, bin[2], bin[1], n_364);
  nand g8 (n_372, n_361, bin[2], bin[1], bin[0]);
  nand g9 (n_373, bin[3], n_362, n_363, n_364);
  nand g10 (n_374, bin[3], n_362, n_363, bin[0]);
  nand g11 (n_375, bin[3], n_362, bin[1], n_364);
  nand g12 (n_376, bin[3], n_362, bin[1], bin[0]);
  nand g13 (n_377, bin[3], bin[2], n_363, n_364);
  nand g14 (n_378, bin[3], bin[2], n_363, bin[0]);
  nand g15 (n_379, bin[3], bin[2], bin[1], n_364);
  nand g16 (n_380, bin[3], bin[2], bin[1], bin[0]);
  not g17 (bitMap[0], n_365);
  not g18 (bitMap[1], n_366);
  not g19 (bitMap[2], n_367);
  not g20 (bitMap[3], n_368);
  not g21 (bitMap[4], n_369);
  not g22 (bitMap[5], n_370);
  not g23 (bitMap[6], n_371);
  not g24 (bitMap[7], n_372);
  not g25 (bitMap[8], n_373);
  not g26 (bitMap[9], n_374);
  not g27 (bitMap[10], n_375);
  not g28 (bitMap[11], n_376);
  not g29 (bitMap[12], n_377);
  not g30 (bitMap[13], n_378);
  not g31 (bitMap[14], n_379);
  not g32 (bitMap[15], n_380);
  not g33 (n_361, bin[3]);
  not g34 (n_362, bin[2]);
  not g35 (n_363, bin[1]);
  not g36 (n_364, bin[0]);
endmodule

module fx68k_or_op(A, Z);
  input [15:0] A;
  output Z;
  wire [15:0] A;
  wire Z;
  wire n_17, n_18, n_19, n_20;
  nor g1 (n_17, A[15], A[14], A[13], A[12]);
  nor g2 (n_18, A[11], A[10], A[9], A[8]);
  nor g3 (n_19, A[7], A[6], A[5], A[4]);
  nor g4 (n_20, A[3], A[2], A[1], A[0]);
  nand g5 (Z, n_17, n_18, n_19, n_20);
endmodule

module fx68k_or_op_4(A, Z);
  input [7:0] A;
  output Z;
  wire [7:0] A;
  wire Z;
  wire n_9, n_10;
  nor g1 (n_10, A[7], A[6], A[5], A[4]);
  nor g2 (n_9, A[3], A[2], A[1], A[0]);
  nand g3 (Z, n_9, n_10);
endmodule

module fx68k_or_op_5(A, Z);
  input [7:0] A;
  output Z;
  wire [7:0] A;
  wire Z;
  wire n_9, n_10;
  nor g1 (n_10, A[7], A[6], A[5], A[4]);
  nor g2 (n_9, A[3], A[2], A[1], A[0]);
  nand g3 (Z, n_9, n_10);
endmodule

module fx68k_case_box_16(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_41(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, z);
  input [8:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  output [9:0] z;
  wire [8:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  wire [9:0] z;
  CDN_mux9 g1(.sel0 (ctl[8]), .data0 (in_0[9]), .sel1 (ctl[7]), .data1
       (in_1[9]), .sel2 (ctl[6]), .data2 (in_2[9]), .sel3 (ctl[5]),
       .data3 (in_3[9]), .sel4 (ctl[4]), .data4 (in_4[9]), .sel5
       (ctl[3]), .data5 (in_5[9]), .sel6 (ctl[2]), .data6 (in_6[9]),
       .sel7 (ctl[1]), .data7 (in_7[9]), .sel8 (ctl[0]), .data8
       (in_8[9]), .z (z[9]));
  CDN_mux9 g11(.sel0 (ctl[8]), .data0 (in_0[8]), .sel1 (ctl[7]), .data1
       (in_1[8]), .sel2 (ctl[6]), .data2 (in_2[8]), .sel3 (ctl[5]),
       .data3 (in_3[8]), .sel4 (ctl[4]), .data4 (in_4[8]), .sel5
       (ctl[3]), .data5 (in_5[8]), .sel6 (ctl[2]), .data6 (in_6[8]),
       .sel7 (ctl[1]), .data7 (in_7[8]), .sel8 (ctl[0]), .data8
       (in_8[8]), .z (z[8]));
  CDN_mux9 g12(.sel0 (ctl[8]), .data0 (in_0[7]), .sel1 (ctl[7]), .data1
       (in_1[7]), .sel2 (ctl[6]), .data2 (in_2[7]), .sel3 (ctl[5]),
       .data3 (in_3[7]), .sel4 (ctl[4]), .data4 (in_4[7]), .sel5
       (ctl[3]), .data5 (in_5[7]), .sel6 (ctl[2]), .data6 (in_6[7]),
       .sel7 (ctl[1]), .data7 (in_7[7]), .sel8 (ctl[0]), .data8
       (in_8[7]), .z (z[7]));
  CDN_mux9 g13(.sel0 (ctl[8]), .data0 (in_0[6]), .sel1 (ctl[7]), .data1
       (in_1[6]), .sel2 (ctl[6]), .data2 (in_2[6]), .sel3 (ctl[5]),
       .data3 (in_3[6]), .sel4 (ctl[4]), .data4 (in_4[6]), .sel5
       (ctl[3]), .data5 (in_5[6]), .sel6 (ctl[2]), .data6 (in_6[6]),
       .sel7 (ctl[1]), .data7 (in_7[6]), .sel8 (ctl[0]), .data8
       (in_8[6]), .z (z[6]));
  CDN_mux9 g14(.sel0 (ctl[8]), .data0 (in_0[5]), .sel1 (ctl[7]), .data1
       (in_1[5]), .sel2 (ctl[6]), .data2 (in_2[5]), .sel3 (ctl[5]),
       .data3 (in_3[5]), .sel4 (ctl[4]), .data4 (in_4[5]), .sel5
       (ctl[3]), .data5 (in_5[5]), .sel6 (ctl[2]), .data6 (in_6[5]),
       .sel7 (ctl[1]), .data7 (in_7[5]), .sel8 (ctl[0]), .data8
       (in_8[5]), .z (z[5]));
  CDN_mux9 g15(.sel0 (ctl[8]), .data0 (in_0[4]), .sel1 (ctl[7]), .data1
       (in_1[4]), .sel2 (ctl[6]), .data2 (in_2[4]), .sel3 (ctl[5]),
       .data3 (in_3[4]), .sel4 (ctl[4]), .data4 (in_4[4]), .sel5
       (ctl[3]), .data5 (in_5[4]), .sel6 (ctl[2]), .data6 (in_6[4]),
       .sel7 (ctl[1]), .data7 (in_7[4]), .sel8 (ctl[0]), .data8
       (in_8[4]), .z (z[4]));
  CDN_mux9 g16(.sel0 (ctl[8]), .data0 (in_0[3]), .sel1 (ctl[7]), .data1
       (in_1[3]), .sel2 (ctl[6]), .data2 (in_2[3]), .sel3 (ctl[5]),
       .data3 (in_3[3]), .sel4 (ctl[4]), .data4 (in_4[3]), .sel5
       (ctl[3]), .data5 (in_5[3]), .sel6 (ctl[2]), .data6 (in_6[3]),
       .sel7 (ctl[1]), .data7 (in_7[3]), .sel8 (ctl[0]), .data8
       (in_8[3]), .z (z[3]));
  CDN_mux9 g17(.sel0 (ctl[8]), .data0 (in_0[2]), .sel1 (ctl[7]), .data1
       (in_1[2]), .sel2 (ctl[6]), .data2 (in_2[2]), .sel3 (ctl[5]),
       .data3 (in_3[2]), .sel4 (ctl[4]), .data4 (in_4[2]), .sel5
       (ctl[3]), .data5 (in_5[2]), .sel6 (ctl[2]), .data6 (in_6[2]),
       .sel7 (ctl[1]), .data7 (in_7[2]), .sel8 (ctl[0]), .data8
       (in_8[2]), .z (z[2]));
  CDN_mux9 g18(.sel0 (ctl[8]), .data0 (in_0[1]), .sel1 (ctl[7]), .data1
       (in_1[1]), .sel2 (ctl[6]), .data2 (in_2[1]), .sel3 (ctl[5]),
       .data3 (in_3[1]), .sel4 (ctl[4]), .data4 (in_4[1]), .sel5
       (ctl[3]), .data5 (in_5[1]), .sel6 (ctl[2]), .data6 (in_6[1]),
       .sel7 (ctl[1]), .data7 (in_7[1]), .sel8 (ctl[0]), .data8
       (in_8[1]), .z (z[1]));
  CDN_mux9 g19(.sel0 (ctl[8]), .data0 (in_0[0]), .sel1 (ctl[7]), .data1
       (in_1[0]), .sel2 (ctl[6]), .data2 (in_2[0]), .sel3 (ctl[5]),
       .data3 (in_3[0]), .sel4 (ctl[4]), .data4 (in_4[0]), .sel5
       (ctl[3]), .data5 (in_5[0]), .sel6 (ctl[2]), .data6 (in_6[0]),
       .sel7 (ctl[1]), .data7 (in_7[0]), .sel8 (ctl[0]), .data8
       (in_8[0]), .z (z[0]));
endmodule

module fx68k_case_box_17(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_20(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_23(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_26(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_77(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [8:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [8:0] z;
  wire [7:0] ctl;
  wire [8:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [8:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[8]), .sel1 (ctl[6]), .data1
       (in_1[8]), .sel2 (ctl[5]), .data2 (in_2[8]), .sel3 (ctl[4]),
       .data3 (in_3[8]), .sel4 (ctl[3]), .data4 (in_4[8]), .sel5
       (ctl[2]), .data5 (in_5[8]), .sel6 (ctl[1]), .data6 (in_6[8]),
       .sel7 (ctl[0]), .data7 (in_7[8]), .z (z[8]));
  CDN_mux8 g10(.sel0 (ctl[7]), .data0 (in_0[7]), .sel1 (ctl[6]), .data1
       (in_1[7]), .sel2 (ctl[5]), .data2 (in_2[7]), .sel3 (ctl[4]),
       .data3 (in_3[7]), .sel4 (ctl[3]), .data4 (in_4[7]), .sel5
       (ctl[2]), .data5 (in_5[7]), .sel6 (ctl[1]), .data6 (in_6[7]),
       .sel7 (ctl[0]), .data7 (in_7[7]), .z (z[7]));
  CDN_mux8 g11(.sel0 (ctl[7]), .data0 (in_0[6]), .sel1 (ctl[6]), .data1
       (in_1[6]), .sel2 (ctl[5]), .data2 (in_2[6]), .sel3 (ctl[4]),
       .data3 (in_3[6]), .sel4 (ctl[3]), .data4 (in_4[6]), .sel5
       (ctl[2]), .data5 (in_5[6]), .sel6 (ctl[1]), .data6 (in_6[6]),
       .sel7 (ctl[0]), .data7 (in_7[6]), .z (z[6]));
  CDN_mux8 g12(.sel0 (ctl[7]), .data0 (in_0[5]), .sel1 (ctl[6]), .data1
       (in_1[5]), .sel2 (ctl[5]), .data2 (in_2[5]), .sel3 (ctl[4]),
       .data3 (in_3[5]), .sel4 (ctl[3]), .data4 (in_4[5]), .sel5
       (ctl[2]), .data5 (in_5[5]), .sel6 (ctl[1]), .data6 (in_6[5]),
       .sel7 (ctl[0]), .data7 (in_7[5]), .z (z[5]));
  CDN_mux8 g13(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g14(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g15(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g16(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g17(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_29(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_32(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_93(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [9:0] z;
  wire [7:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [9:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[9]), .sel1 (ctl[6]), .data1
       (in_1[9]), .sel2 (ctl[5]), .data2 (in_2[9]), .sel3 (ctl[4]),
       .data3 (in_3[9]), .sel4 (ctl[3]), .data4 (in_4[9]), .sel5
       (ctl[2]), .data5 (in_5[9]), .sel6 (ctl[1]), .data6 (in_6[9]),
       .sel7 (ctl[0]), .data7 (in_7[9]), .z (z[9]));
  CDN_mux8 g11(.sel0 (ctl[7]), .data0 (in_0[8]), .sel1 (ctl[6]), .data1
       (in_1[8]), .sel2 (ctl[5]), .data2 (in_2[8]), .sel3 (ctl[4]),
       .data3 (in_3[8]), .sel4 (ctl[3]), .data4 (in_4[8]), .sel5
       (ctl[2]), .data5 (in_5[8]), .sel6 (ctl[1]), .data6 (in_6[8]),
       .sel7 (ctl[0]), .data7 (in_7[8]), .z (z[8]));
  CDN_mux8 g12(.sel0 (ctl[7]), .data0 (in_0[7]), .sel1 (ctl[6]), .data1
       (in_1[7]), .sel2 (ctl[5]), .data2 (in_2[7]), .sel3 (ctl[4]),
       .data3 (in_3[7]), .sel4 (ctl[3]), .data4 (in_4[7]), .sel5
       (ctl[2]), .data5 (in_5[7]), .sel6 (ctl[1]), .data6 (in_6[7]),
       .sel7 (ctl[0]), .data7 (in_7[7]), .z (z[7]));
  CDN_mux8 g13(.sel0 (ctl[7]), .data0 (in_0[6]), .sel1 (ctl[6]), .data1
       (in_1[6]), .sel2 (ctl[5]), .data2 (in_2[6]), .sel3 (ctl[4]),
       .data3 (in_3[6]), .sel4 (ctl[3]), .data4 (in_4[6]), .sel5
       (ctl[2]), .data5 (in_5[6]), .sel6 (ctl[1]), .data6 (in_6[6]),
       .sel7 (ctl[0]), .data7 (in_7[6]), .z (z[6]));
  CDN_mux8 g14(.sel0 (ctl[7]), .data0 (in_0[5]), .sel1 (ctl[6]), .data1
       (in_1[5]), .sel2 (ctl[5]), .data2 (in_2[5]), .sel3 (ctl[4]),
       .data3 (in_3[5]), .sel4 (ctl[3]), .data4 (in_4[5]), .sel5
       (ctl[2]), .data5 (in_5[5]), .sel6 (ctl[1]), .data6 (in_6[5]),
       .sel7 (ctl[0]), .data7 (in_7[5]), .z (z[5]));
  CDN_mux8 g15(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g16(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g17(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g18(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g19(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_35(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_38(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_41(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_119(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  output [9:0] z;
  wire [11:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  wire [9:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[9]), .sel1 (ctl[10]),
       .data1 (in_1[9]), .sel2 (ctl[9]), .data2 (in_2[9]), .sel3
       (ctl[8]), .data3 (in_3[9]), .sel4 (ctl[7]), .data4 (in_4[9]),
       .sel5 (ctl[6]), .data5 (in_5[9]), .sel6 (ctl[5]), .data6
       (in_6[9]), .sel7 (ctl[4]), .data7 (in_7[9]), .sel8 (ctl[3]),
       .data8 (in_8[9]), .sel9 (ctl[2]), .data9 (in_9[9]), .sel10
       (ctl[1]), .data10 (in_10[9]), .sel11 (ctl[0]), .data11
       (in_11[9]), .z (z[9]));
  CDN_mux12 g11(.sel0 (ctl[11]), .data0 (in_0[8]), .sel1 (ctl[10]),
       .data1 (in_1[8]), .sel2 (ctl[9]), .data2 (in_2[8]), .sel3
       (ctl[8]), .data3 (in_3[8]), .sel4 (ctl[7]), .data4 (in_4[8]),
       .sel5 (ctl[6]), .data5 (in_5[8]), .sel6 (ctl[5]), .data6
       (in_6[8]), .sel7 (ctl[4]), .data7 (in_7[8]), .sel8 (ctl[3]),
       .data8 (in_8[8]), .sel9 (ctl[2]), .data9 (in_9[8]), .sel10
       (ctl[1]), .data10 (in_10[8]), .sel11 (ctl[0]), .data11
       (in_11[8]), .z (z[8]));
  CDN_mux12 g12(.sel0 (ctl[11]), .data0 (in_0[7]), .sel1 (ctl[10]),
       .data1 (in_1[7]), .sel2 (ctl[9]), .data2 (in_2[7]), .sel3
       (ctl[8]), .data3 (in_3[7]), .sel4 (ctl[7]), .data4 (in_4[7]),
       .sel5 (ctl[6]), .data5 (in_5[7]), .sel6 (ctl[5]), .data6
       (in_6[7]), .sel7 (ctl[4]), .data7 (in_7[7]), .sel8 (ctl[3]),
       .data8 (in_8[7]), .sel9 (ctl[2]), .data9 (in_9[7]), .sel10
       (ctl[1]), .data10 (in_10[7]), .sel11 (ctl[0]), .data11
       (in_11[7]), .z (z[7]));
  CDN_mux12 g13(.sel0 (ctl[11]), .data0 (in_0[6]), .sel1 (ctl[10]),
       .data1 (in_1[6]), .sel2 (ctl[9]), .data2 (in_2[6]), .sel3
       (ctl[8]), .data3 (in_3[6]), .sel4 (ctl[7]), .data4 (in_4[6]),
       .sel5 (ctl[6]), .data5 (in_5[6]), .sel6 (ctl[5]), .data6
       (in_6[6]), .sel7 (ctl[4]), .data7 (in_7[6]), .sel8 (ctl[3]),
       .data8 (in_8[6]), .sel9 (ctl[2]), .data9 (in_9[6]), .sel10
       (ctl[1]), .data10 (in_10[6]), .sel11 (ctl[0]), .data11
       (in_11[6]), .z (z[6]));
  CDN_mux12 g14(.sel0 (ctl[11]), .data0 (in_0[5]), .sel1 (ctl[10]),
       .data1 (in_1[5]), .sel2 (ctl[9]), .data2 (in_2[5]), .sel3
       (ctl[8]), .data3 (in_3[5]), .sel4 (ctl[7]), .data4 (in_4[5]),
       .sel5 (ctl[6]), .data5 (in_5[5]), .sel6 (ctl[5]), .data6
       (in_6[5]), .sel7 (ctl[4]), .data7 (in_7[5]), .sel8 (ctl[3]),
       .data8 (in_8[5]), .sel9 (ctl[2]), .data9 (in_9[5]), .sel10
       (ctl[1]), .data10 (in_10[5]), .sel11 (ctl[0]), .data11
       (in_11[5]), .z (z[5]));
  CDN_mux12 g15(.sel0 (ctl[11]), .data0 (in_0[4]), .sel1 (ctl[10]),
       .data1 (in_1[4]), .sel2 (ctl[9]), .data2 (in_2[4]), .sel3
       (ctl[8]), .data3 (in_3[4]), .sel4 (ctl[7]), .data4 (in_4[4]),
       .sel5 (ctl[6]), .data5 (in_5[4]), .sel6 (ctl[5]), .data6
       (in_6[4]), .sel7 (ctl[4]), .data7 (in_7[4]), .sel8 (ctl[3]),
       .data8 (in_8[4]), .sel9 (ctl[2]), .data9 (in_9[4]), .sel10
       (ctl[1]), .data10 (in_10[4]), .sel11 (ctl[0]), .data11
       (in_11[4]), .z (z[4]));
  CDN_mux12 g16(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g17(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g18(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g19(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_case_box_44(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_128(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, z);
  input [8:0] ctl;
  input [19:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  output [19:0] z;
  wire [8:0] ctl;
  wire [19:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  wire [19:0] z;
  CDN_mux9 g1(.sel0 (ctl[8]), .data0 (in_0[19]), .sel1 (ctl[7]), .data1
       (in_1[19]), .sel2 (ctl[6]), .data2 (in_2[19]), .sel3 (ctl[5]),
       .data3 (in_3[19]), .sel4 (ctl[4]), .data4 (in_4[19]), .sel5
       (ctl[3]), .data5 (in_5[19]), .sel6 (ctl[2]), .data6 (in_6[19]),
       .sel7 (ctl[1]), .data7 (in_7[19]), .sel8 (ctl[0]), .data8
       (in_8[19]), .z (z[19]));
  CDN_mux9 g21(.sel0 (ctl[8]), .data0 (in_0[18]), .sel1 (ctl[7]),
       .data1 (in_1[18]), .sel2 (ctl[6]), .data2 (in_2[18]), .sel3
       (ctl[5]), .data3 (in_3[18]), .sel4 (ctl[4]), .data4 (in_4[18]),
       .sel5 (ctl[3]), .data5 (in_5[18]), .sel6 (ctl[2]), .data6
       (in_6[18]), .sel7 (ctl[1]), .data7 (in_7[18]), .sel8 (ctl[0]),
       .data8 (in_8[18]), .z (z[18]));
  CDN_mux9 g22(.sel0 (ctl[8]), .data0 (in_0[17]), .sel1 (ctl[7]),
       .data1 (in_1[17]), .sel2 (ctl[6]), .data2 (in_2[17]), .sel3
       (ctl[5]), .data3 (in_3[17]), .sel4 (ctl[4]), .data4 (in_4[17]),
       .sel5 (ctl[3]), .data5 (in_5[17]), .sel6 (ctl[2]), .data6
       (in_6[17]), .sel7 (ctl[1]), .data7 (in_7[17]), .sel8 (ctl[0]),
       .data8 (in_8[17]), .z (z[17]));
  CDN_mux9 g23(.sel0 (ctl[8]), .data0 (in_0[16]), .sel1 (ctl[7]),
       .data1 (in_1[16]), .sel2 (ctl[6]), .data2 (in_2[16]), .sel3
       (ctl[5]), .data3 (in_3[16]), .sel4 (ctl[4]), .data4 (in_4[16]),
       .sel5 (ctl[3]), .data5 (in_5[16]), .sel6 (ctl[2]), .data6
       (in_6[16]), .sel7 (ctl[1]), .data7 (in_7[16]), .sel8 (ctl[0]),
       .data8 (in_8[16]), .z (z[16]));
  CDN_mux9 g24(.sel0 (ctl[8]), .data0 (in_0[15]), .sel1 (ctl[7]),
       .data1 (in_1[15]), .sel2 (ctl[6]), .data2 (in_2[15]), .sel3
       (ctl[5]), .data3 (in_3[15]), .sel4 (ctl[4]), .data4 (in_4[15]),
       .sel5 (ctl[3]), .data5 (in_5[15]), .sel6 (ctl[2]), .data6
       (in_6[15]), .sel7 (ctl[1]), .data7 (in_7[15]), .sel8 (ctl[0]),
       .data8 (in_8[15]), .z (z[15]));
  CDN_mux9 g25(.sel0 (ctl[8]), .data0 (in_0[14]), .sel1 (ctl[7]),
       .data1 (in_1[14]), .sel2 (ctl[6]), .data2 (in_2[14]), .sel3
       (ctl[5]), .data3 (in_3[14]), .sel4 (ctl[4]), .data4 (in_4[14]),
       .sel5 (ctl[3]), .data5 (in_5[14]), .sel6 (ctl[2]), .data6
       (in_6[14]), .sel7 (ctl[1]), .data7 (in_7[14]), .sel8 (ctl[0]),
       .data8 (in_8[14]), .z (z[14]));
  CDN_mux9 g26(.sel0 (ctl[8]), .data0 (in_0[13]), .sel1 (ctl[7]),
       .data1 (in_1[13]), .sel2 (ctl[6]), .data2 (in_2[13]), .sel3
       (ctl[5]), .data3 (in_3[13]), .sel4 (ctl[4]), .data4 (in_4[13]),
       .sel5 (ctl[3]), .data5 (in_5[13]), .sel6 (ctl[2]), .data6
       (in_6[13]), .sel7 (ctl[1]), .data7 (in_7[13]), .sel8 (ctl[0]),
       .data8 (in_8[13]), .z (z[13]));
  CDN_mux9 g27(.sel0 (ctl[8]), .data0 (in_0[12]), .sel1 (ctl[7]),
       .data1 (in_1[12]), .sel2 (ctl[6]), .data2 (in_2[12]), .sel3
       (ctl[5]), .data3 (in_3[12]), .sel4 (ctl[4]), .data4 (in_4[12]),
       .sel5 (ctl[3]), .data5 (in_5[12]), .sel6 (ctl[2]), .data6
       (in_6[12]), .sel7 (ctl[1]), .data7 (in_7[12]), .sel8 (ctl[0]),
       .data8 (in_8[12]), .z (z[12]));
  CDN_mux9 g28(.sel0 (ctl[8]), .data0 (in_0[11]), .sel1 (ctl[7]),
       .data1 (in_1[11]), .sel2 (ctl[6]), .data2 (in_2[11]), .sel3
       (ctl[5]), .data3 (in_3[11]), .sel4 (ctl[4]), .data4 (in_4[11]),
       .sel5 (ctl[3]), .data5 (in_5[11]), .sel6 (ctl[2]), .data6
       (in_6[11]), .sel7 (ctl[1]), .data7 (in_7[11]), .sel8 (ctl[0]),
       .data8 (in_8[11]), .z (z[11]));
  CDN_mux9 g29(.sel0 (ctl[8]), .data0 (in_0[10]), .sel1 (ctl[7]),
       .data1 (in_1[10]), .sel2 (ctl[6]), .data2 (in_2[10]), .sel3
       (ctl[5]), .data3 (in_3[10]), .sel4 (ctl[4]), .data4 (in_4[10]),
       .sel5 (ctl[3]), .data5 (in_5[10]), .sel6 (ctl[2]), .data6
       (in_6[10]), .sel7 (ctl[1]), .data7 (in_7[10]), .sel8 (ctl[0]),
       .data8 (in_8[10]), .z (z[10]));
  CDN_mux9 g30(.sel0 (ctl[8]), .data0 (in_0[9]), .sel1 (ctl[7]), .data1
       (in_1[9]), .sel2 (ctl[6]), .data2 (in_2[9]), .sel3 (ctl[5]),
       .data3 (in_3[9]), .sel4 (ctl[4]), .data4 (in_4[9]), .sel5
       (ctl[3]), .data5 (in_5[9]), .sel6 (ctl[2]), .data6 (in_6[9]),
       .sel7 (ctl[1]), .data7 (in_7[9]), .sel8 (ctl[0]), .data8
       (in_8[9]), .z (z[9]));
  CDN_mux9 g31(.sel0 (ctl[8]), .data0 (in_0[8]), .sel1 (ctl[7]), .data1
       (in_1[8]), .sel2 (ctl[6]), .data2 (in_2[8]), .sel3 (ctl[5]),
       .data3 (in_3[8]), .sel4 (ctl[4]), .data4 (in_4[8]), .sel5
       (ctl[3]), .data5 (in_5[8]), .sel6 (ctl[2]), .data6 (in_6[8]),
       .sel7 (ctl[1]), .data7 (in_7[8]), .sel8 (ctl[0]), .data8
       (in_8[8]), .z (z[8]));
  CDN_mux9 g32(.sel0 (ctl[8]), .data0 (in_0[7]), .sel1 (ctl[7]), .data1
       (in_1[7]), .sel2 (ctl[6]), .data2 (in_2[7]), .sel3 (ctl[5]),
       .data3 (in_3[7]), .sel4 (ctl[4]), .data4 (in_4[7]), .sel5
       (ctl[3]), .data5 (in_5[7]), .sel6 (ctl[2]), .data6 (in_6[7]),
       .sel7 (ctl[1]), .data7 (in_7[7]), .sel8 (ctl[0]), .data8
       (in_8[7]), .z (z[7]));
  CDN_mux9 g33(.sel0 (ctl[8]), .data0 (in_0[6]), .sel1 (ctl[7]), .data1
       (in_1[6]), .sel2 (ctl[6]), .data2 (in_2[6]), .sel3 (ctl[5]),
       .data3 (in_3[6]), .sel4 (ctl[4]), .data4 (in_4[6]), .sel5
       (ctl[3]), .data5 (in_5[6]), .sel6 (ctl[2]), .data6 (in_6[6]),
       .sel7 (ctl[1]), .data7 (in_7[6]), .sel8 (ctl[0]), .data8
       (in_8[6]), .z (z[6]));
  CDN_mux9 g34(.sel0 (ctl[8]), .data0 (in_0[5]), .sel1 (ctl[7]), .data1
       (in_1[5]), .sel2 (ctl[6]), .data2 (in_2[5]), .sel3 (ctl[5]),
       .data3 (in_3[5]), .sel4 (ctl[4]), .data4 (in_4[5]), .sel5
       (ctl[3]), .data5 (in_5[5]), .sel6 (ctl[2]), .data6 (in_6[5]),
       .sel7 (ctl[1]), .data7 (in_7[5]), .sel8 (ctl[0]), .data8
       (in_8[5]), .z (z[5]));
  CDN_mux9 g35(.sel0 (ctl[8]), .data0 (in_0[4]), .sel1 (ctl[7]), .data1
       (in_1[4]), .sel2 (ctl[6]), .data2 (in_2[4]), .sel3 (ctl[5]),
       .data3 (in_3[4]), .sel4 (ctl[4]), .data4 (in_4[4]), .sel5
       (ctl[3]), .data5 (in_5[4]), .sel6 (ctl[2]), .data6 (in_6[4]),
       .sel7 (ctl[1]), .data7 (in_7[4]), .sel8 (ctl[0]), .data8
       (in_8[4]), .z (z[4]));
  CDN_mux9 g36(.sel0 (ctl[8]), .data0 (in_0[3]), .sel1 (ctl[7]), .data1
       (in_1[3]), .sel2 (ctl[6]), .data2 (in_2[3]), .sel3 (ctl[5]),
       .data3 (in_3[3]), .sel4 (ctl[4]), .data4 (in_4[3]), .sel5
       (ctl[3]), .data5 (in_5[3]), .sel6 (ctl[2]), .data6 (in_6[3]),
       .sel7 (ctl[1]), .data7 (in_7[3]), .sel8 (ctl[0]), .data8
       (in_8[3]), .z (z[3]));
  CDN_mux9 g37(.sel0 (ctl[8]), .data0 (in_0[2]), .sel1 (ctl[7]), .data1
       (in_1[2]), .sel2 (ctl[6]), .data2 (in_2[2]), .sel3 (ctl[5]),
       .data3 (in_3[2]), .sel4 (ctl[4]), .data4 (in_4[2]), .sel5
       (ctl[3]), .data5 (in_5[2]), .sel6 (ctl[2]), .data6 (in_6[2]),
       .sel7 (ctl[1]), .data7 (in_7[2]), .sel8 (ctl[0]), .data8
       (in_8[2]), .z (z[2]));
  CDN_mux9 g38(.sel0 (ctl[8]), .data0 (in_0[1]), .sel1 (ctl[7]), .data1
       (in_1[1]), .sel2 (ctl[6]), .data2 (in_2[1]), .sel3 (ctl[5]),
       .data3 (in_3[1]), .sel4 (ctl[4]), .data4 (in_4[1]), .sel5
       (ctl[3]), .data5 (in_5[1]), .sel6 (ctl[2]), .data6 (in_6[1]),
       .sel7 (ctl[1]), .data7 (in_7[1]), .sel8 (ctl[0]), .data8
       (in_8[1]), .z (z[1]));
  CDN_mux9 g39(.sel0 (ctl[8]), .data0 (in_0[0]), .sel1 (ctl[7]), .data1
       (in_1[0]), .sel2 (ctl[6]), .data2 (in_2[0]), .sel3 (ctl[5]),
       .data3 (in_3[0]), .sel4 (ctl[4]), .data4 (in_4[0]), .sel5
       (ctl[3]), .data5 (in_5[0]), .sel6 (ctl[2]), .data6 (in_6[0]),
       .sel7 (ctl[1]), .data7 (in_7[0]), .sel8 (ctl[0]), .data8
       (in_8[0]), .z (z[0]));
endmodule

module fx68k_case_box_47(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_50(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_53(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_185(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, z);
  input [9:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7,
       in_8, in_9;
  output [9:0] z;
  wire [9:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9;
  wire [9:0] z;
  CDN_mux10 g1(.sel0 (ctl[9]), .data0 (in_0[9]), .sel1 (ctl[8]), .data1
       (in_1[9]), .sel2 (ctl[7]), .data2 (in_2[9]), .sel3 (ctl[6]),
       .data3 (in_3[9]), .sel4 (ctl[5]), .data4 (in_4[9]), .sel5
       (ctl[4]), .data5 (in_5[9]), .sel6 (ctl[3]), .data6 (in_6[9]),
       .sel7 (ctl[2]), .data7 (in_7[9]), .sel8 (ctl[1]), .data8
       (in_8[9]), .sel9 (ctl[0]), .data9 (in_9[9]), .z (z[9]));
  CDN_mux10 g11(.sel0 (ctl[9]), .data0 (in_0[8]), .sel1 (ctl[8]),
       .data1 (in_1[8]), .sel2 (ctl[7]), .data2 (in_2[8]), .sel3
       (ctl[6]), .data3 (in_3[8]), .sel4 (ctl[5]), .data4 (in_4[8]),
       .sel5 (ctl[4]), .data5 (in_5[8]), .sel6 (ctl[3]), .data6
       (in_6[8]), .sel7 (ctl[2]), .data7 (in_7[8]), .sel8 (ctl[1]),
       .data8 (in_8[8]), .sel9 (ctl[0]), .data9 (in_9[8]), .z (z[8]));
  CDN_mux10 g12(.sel0 (ctl[9]), .data0 (in_0[7]), .sel1 (ctl[8]),
       .data1 (in_1[7]), .sel2 (ctl[7]), .data2 (in_2[7]), .sel3
       (ctl[6]), .data3 (in_3[7]), .sel4 (ctl[5]), .data4 (in_4[7]),
       .sel5 (ctl[4]), .data5 (in_5[7]), .sel6 (ctl[3]), .data6
       (in_6[7]), .sel7 (ctl[2]), .data7 (in_7[7]), .sel8 (ctl[1]),
       .data8 (in_8[7]), .sel9 (ctl[0]), .data9 (in_9[7]), .z (z[7]));
  CDN_mux10 g13(.sel0 (ctl[9]), .data0 (in_0[6]), .sel1 (ctl[8]),
       .data1 (in_1[6]), .sel2 (ctl[7]), .data2 (in_2[6]), .sel3
       (ctl[6]), .data3 (in_3[6]), .sel4 (ctl[5]), .data4 (in_4[6]),
       .sel5 (ctl[4]), .data5 (in_5[6]), .sel6 (ctl[3]), .data6
       (in_6[6]), .sel7 (ctl[2]), .data7 (in_7[6]), .sel8 (ctl[1]),
       .data8 (in_8[6]), .sel9 (ctl[0]), .data9 (in_9[6]), .z (z[6]));
  CDN_mux10 g14(.sel0 (ctl[9]), .data0 (in_0[5]), .sel1 (ctl[8]),
       .data1 (in_1[5]), .sel2 (ctl[7]), .data2 (in_2[5]), .sel3
       (ctl[6]), .data3 (in_3[5]), .sel4 (ctl[5]), .data4 (in_4[5]),
       .sel5 (ctl[4]), .data5 (in_5[5]), .sel6 (ctl[3]), .data6
       (in_6[5]), .sel7 (ctl[2]), .data7 (in_7[5]), .sel8 (ctl[1]),
       .data8 (in_8[5]), .sel9 (ctl[0]), .data9 (in_9[5]), .z (z[5]));
  CDN_mux10 g15(.sel0 (ctl[9]), .data0 (in_0[4]), .sel1 (ctl[8]),
       .data1 (in_1[4]), .sel2 (ctl[7]), .data2 (in_2[4]), .sel3
       (ctl[6]), .data3 (in_3[4]), .sel4 (ctl[5]), .data4 (in_4[4]),
       .sel5 (ctl[4]), .data5 (in_5[4]), .sel6 (ctl[3]), .data6
       (in_6[4]), .sel7 (ctl[2]), .data7 (in_7[4]), .sel8 (ctl[1]),
       .data8 (in_8[4]), .sel9 (ctl[0]), .data9 (in_9[4]), .z (z[4]));
  CDN_mux10 g16(.sel0 (ctl[9]), .data0 (in_0[3]), .sel1 (ctl[8]),
       .data1 (in_1[3]), .sel2 (ctl[7]), .data2 (in_2[3]), .sel3
       (ctl[6]), .data3 (in_3[3]), .sel4 (ctl[5]), .data4 (in_4[3]),
       .sel5 (ctl[4]), .data5 (in_5[3]), .sel6 (ctl[3]), .data6
       (in_6[3]), .sel7 (ctl[2]), .data7 (in_7[3]), .sel8 (ctl[1]),
       .data8 (in_8[3]), .sel9 (ctl[0]), .data9 (in_9[3]), .z (z[3]));
  CDN_mux10 g17(.sel0 (ctl[9]), .data0 (in_0[2]), .sel1 (ctl[8]),
       .data1 (in_1[2]), .sel2 (ctl[7]), .data2 (in_2[2]), .sel3
       (ctl[6]), .data3 (in_3[2]), .sel4 (ctl[5]), .data4 (in_4[2]),
       .sel5 (ctl[4]), .data5 (in_5[2]), .sel6 (ctl[3]), .data6
       (in_6[2]), .sel7 (ctl[2]), .data7 (in_7[2]), .sel8 (ctl[1]),
       .data8 (in_8[2]), .sel9 (ctl[0]), .data9 (in_9[2]), .z (z[2]));
  CDN_mux10 g18(.sel0 (ctl[9]), .data0 (in_0[1]), .sel1 (ctl[8]),
       .data1 (in_1[1]), .sel2 (ctl[7]), .data2 (in_2[1]), .sel3
       (ctl[6]), .data3 (in_3[1]), .sel4 (ctl[5]), .data4 (in_4[1]),
       .sel5 (ctl[4]), .data5 (in_5[1]), .sel6 (ctl[3]), .data6
       (in_6[1]), .sel7 (ctl[2]), .data7 (in_7[1]), .sel8 (ctl[1]),
       .data8 (in_8[1]), .sel9 (ctl[0]), .data9 (in_9[1]), .z (z[1]));
  CDN_mux10 g19(.sel0 (ctl[9]), .data0 (in_0[0]), .sel1 (ctl[8]),
       .data1 (in_1[0]), .sel2 (ctl[7]), .data2 (in_2[0]), .sel3
       (ctl[6]), .data3 (in_3[0]), .sel4 (ctl[5]), .data4 (in_4[0]),
       .sel5 (ctl[4]), .data5 (in_5[0]), .sel6 (ctl[3]), .data6
       (in_6[0]), .sel7 (ctl[2]), .data7 (in_7[0]), .sel8 (ctl[1]),
       .data8 (in_8[0]), .sel9 (ctl[0]), .data9 (in_9[0]), .z (z[0]));
endmodule

module fx68k_case_box_56(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_59(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_62(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_65(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_68(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_71(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_247(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [7:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [7:0] z;
  wire [6:0] ctl;
  wire [7:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [7:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[7]), .sel1 (ctl[5]), .data1
       (in_1[7]), .sel2 (ctl[4]), .data2 (in_2[7]), .sel3 (ctl[3]),
       .data3 (in_3[7]), .sel4 (ctl[2]), .data4 (in_4[7]), .sel5
       (ctl[1]), .data5 (in_5[7]), .sel6 (ctl[0]), .data6 (in_6[7]), .z
       (z[7]));
  CDN_mux7 g9(.sel0 (ctl[6]), .data0 (in_0[6]), .sel1 (ctl[5]), .data1
       (in_1[6]), .sel2 (ctl[4]), .data2 (in_2[6]), .sel3 (ctl[3]),
       .data3 (in_3[6]), .sel4 (ctl[2]), .data4 (in_4[6]), .sel5
       (ctl[1]), .data5 (in_5[6]), .sel6 (ctl[0]), .data6 (in_6[6]), .z
       (z[6]));
  CDN_mux7 g10(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g11(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g12(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g13(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g14(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g15(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_mux_254(ctl, in_0, in_1, in_2, in_3, in_4, z);
  input [4:0] ctl;
  input [7:0] in_0, in_1, in_2, in_3, in_4;
  output [7:0] z;
  wire [4:0] ctl;
  wire [7:0] in_0, in_1, in_2, in_3, in_4;
  wire [7:0] z;
  CDN_mux5 g1(.sel0 (ctl[4]), .data0 (in_0[7]), .sel1 (ctl[3]), .data1
       (in_1[7]), .sel2 (ctl[2]), .data2 (in_2[7]), .sel3 (ctl[1]),
       .data3 (in_3[7]), .sel4 (ctl[0]), .data4 (in_4[7]), .z (z[7]));
  CDN_mux5 g9(.sel0 (ctl[4]), .data0 (in_0[6]), .sel1 (ctl[3]), .data1
       (in_1[6]), .sel2 (ctl[2]), .data2 (in_2[6]), .sel3 (ctl[1]),
       .data3 (in_3[6]), .sel4 (ctl[0]), .data4 (in_4[6]), .z (z[6]));
  CDN_mux5 g10(.sel0 (ctl[4]), .data0 (in_0[5]), .sel1 (ctl[3]), .data1
       (in_1[5]), .sel2 (ctl[2]), .data2 (in_2[5]), .sel3 (ctl[1]),
       .data3 (in_3[5]), .sel4 (ctl[0]), .data4 (in_4[5]), .z (z[5]));
  CDN_mux5 g11(.sel0 (ctl[4]), .data0 (in_0[4]), .sel1 (ctl[3]), .data1
       (in_1[4]), .sel2 (ctl[2]), .data2 (in_2[4]), .sel3 (ctl[1]),
       .data3 (in_3[4]), .sel4 (ctl[0]), .data4 (in_4[4]), .z (z[4]));
  CDN_mux5 g12(.sel0 (ctl[4]), .data0 (in_0[3]), .sel1 (ctl[3]), .data1
       (in_1[3]), .sel2 (ctl[2]), .data2 (in_2[3]), .sel3 (ctl[1]),
       .data3 (in_3[3]), .sel4 (ctl[0]), .data4 (in_4[3]), .z (z[3]));
  CDN_mux5 g13(.sel0 (ctl[4]), .data0 (in_0[2]), .sel1 (ctl[3]), .data1
       (in_1[2]), .sel2 (ctl[2]), .data2 (in_2[2]), .sel3 (ctl[1]),
       .data3 (in_3[2]), .sel4 (ctl[0]), .data4 (in_4[2]), .z (z[2]));
  CDN_mux5 g14(.sel0 (ctl[4]), .data0 (in_0[1]), .sel1 (ctl[3]), .data1
       (in_1[1]), .sel2 (ctl[2]), .data2 (in_2[1]), .sel3 (ctl[1]),
       .data3 (in_3[1]), .sel4 (ctl[0]), .data4 (in_4[1]), .z (z[1]));
  CDN_mux5 g15(.sel0 (ctl[4]), .data0 (in_0[0]), .sel1 (ctl[3]), .data1
       (in_1[0]), .sel2 (ctl[2]), .data2 (in_2[0]), .sel3 (ctl[1]),
       .data3 (in_3[0]), .sel4 (ctl[0]), .data4 (in_4[0]), .z (z[0]));
endmodule

module fx68k_bmux(ctl, in_0, in_1, z);
  input ctl;
  input [7:0] in_0, in_1;
  output [7:0] z;
  wire ctl;
  wire [7:0] in_0, in_1;
  wire [7:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[7]), .data1 (in_1[7]), .z
       (z[7]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[6]), .data1 (in_1[6]), .z
       (z[6]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g7(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g8(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_mux_272(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [9:0] z;
  wire [6:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [9:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[9]), .sel1 (ctl[5]), .data1
       (in_1[9]), .sel2 (ctl[4]), .data2 (in_2[9]), .sel3 (ctl[3]),
       .data3 (in_3[9]), .sel4 (ctl[2]), .data4 (in_4[9]), .sel5
       (ctl[1]), .data5 (in_5[9]), .sel6 (ctl[0]), .data6 (in_6[9]), .z
       (z[9]));
  CDN_mux7 g11(.sel0 (ctl[6]), .data0 (in_0[8]), .sel1 (ctl[5]), .data1
       (in_1[8]), .sel2 (ctl[4]), .data2 (in_2[8]), .sel3 (ctl[3]),
       .data3 (in_3[8]), .sel4 (ctl[2]), .data4 (in_4[8]), .sel5
       (ctl[1]), .data5 (in_5[8]), .sel6 (ctl[0]), .data6 (in_6[8]), .z
       (z[8]));
  CDN_mux7 g12(.sel0 (ctl[6]), .data0 (in_0[7]), .sel1 (ctl[5]), .data1
       (in_1[7]), .sel2 (ctl[4]), .data2 (in_2[7]), .sel3 (ctl[3]),
       .data3 (in_3[7]), .sel4 (ctl[2]), .data4 (in_4[7]), .sel5
       (ctl[1]), .data5 (in_5[7]), .sel6 (ctl[0]), .data6 (in_6[7]), .z
       (z[7]));
  CDN_mux7 g13(.sel0 (ctl[6]), .data0 (in_0[6]), .sel1 (ctl[5]), .data1
       (in_1[6]), .sel2 (ctl[4]), .data2 (in_2[6]), .sel3 (ctl[3]),
       .data3 (in_3[6]), .sel4 (ctl[2]), .data4 (in_4[6]), .sel5
       (ctl[1]), .data5 (in_5[6]), .sel6 (ctl[0]), .data6 (in_6[6]), .z
       (z[6]));
  CDN_mux7 g14(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g15(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g16(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g17(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g18(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g19(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_mux_281(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input [9:0] in_0, in_1;
  output [9:0] z;
  wire [1:0] ctl;
  wire [9:0] in_0, in_1;
  wire [9:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[9]), .sel1 (ctl[0]), .data1
       (in_1[9]), .z (z[9]));
  CDN_mux2 g11(.sel0 (ctl[1]), .data0 (in_0[8]), .sel1 (ctl[0]), .data1
       (in_1[8]), .z (z[8]));
  CDN_mux2 g12(.sel0 (ctl[1]), .data0 (in_0[7]), .sel1 (ctl[0]), .data1
       (in_1[7]), .z (z[7]));
  CDN_mux2 g13(.sel0 (ctl[1]), .data0 (in_0[6]), .sel1 (ctl[0]), .data1
       (in_1[6]), .z (z[6]));
  CDN_mux2 g14(.sel0 (ctl[1]), .data0 (in_0[5]), .sel1 (ctl[0]), .data1
       (in_1[5]), .z (z[5]));
  CDN_mux2 g15(.sel0 (ctl[1]), .data0 (in_0[4]), .sel1 (ctl[0]), .data1
       (in_1[4]), .z (z[4]));
  CDN_mux2 g16(.sel0 (ctl[1]), .data0 (in_0[3]), .sel1 (ctl[0]), .data1
       (in_1[3]), .z (z[3]));
  CDN_mux2 g17(.sel0 (ctl[1]), .data0 (in_0[2]), .sel1 (ctl[0]), .data1
       (in_1[2]), .z (z[2]));
  CDN_mux2 g18(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g19(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_mux_290(ctl, in_0, in_1, in_2, in_3, in_4, z);
  input [4:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4;
  output [9:0] z;
  wire [4:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4;
  wire [9:0] z;
  CDN_mux5 g1(.sel0 (ctl[4]), .data0 (in_0[9]), .sel1 (ctl[3]), .data1
       (in_1[9]), .sel2 (ctl[2]), .data2 (in_2[9]), .sel3 (ctl[1]),
       .data3 (in_3[9]), .sel4 (ctl[0]), .data4 (in_4[9]), .z (z[9]));
  CDN_mux5 g11(.sel0 (ctl[4]), .data0 (in_0[8]), .sel1 (ctl[3]), .data1
       (in_1[8]), .sel2 (ctl[2]), .data2 (in_2[8]), .sel3 (ctl[1]),
       .data3 (in_3[8]), .sel4 (ctl[0]), .data4 (in_4[8]), .z (z[8]));
  CDN_mux5 g12(.sel0 (ctl[4]), .data0 (in_0[7]), .sel1 (ctl[3]), .data1
       (in_1[7]), .sel2 (ctl[2]), .data2 (in_2[7]), .sel3 (ctl[1]),
       .data3 (in_3[7]), .sel4 (ctl[0]), .data4 (in_4[7]), .z (z[7]));
  CDN_mux5 g13(.sel0 (ctl[4]), .data0 (in_0[6]), .sel1 (ctl[3]), .data1
       (in_1[6]), .sel2 (ctl[2]), .data2 (in_2[6]), .sel3 (ctl[1]),
       .data3 (in_3[6]), .sel4 (ctl[0]), .data4 (in_4[6]), .z (z[6]));
  CDN_mux5 g14(.sel0 (ctl[4]), .data0 (in_0[5]), .sel1 (ctl[3]), .data1
       (in_1[5]), .sel2 (ctl[2]), .data2 (in_2[5]), .sel3 (ctl[1]),
       .data3 (in_3[5]), .sel4 (ctl[0]), .data4 (in_4[5]), .z (z[5]));
  CDN_mux5 g15(.sel0 (ctl[4]), .data0 (in_0[4]), .sel1 (ctl[3]), .data1
       (in_1[4]), .sel2 (ctl[2]), .data2 (in_2[4]), .sel3 (ctl[1]),
       .data3 (in_3[4]), .sel4 (ctl[0]), .data4 (in_4[4]), .z (z[4]));
  CDN_mux5 g16(.sel0 (ctl[4]), .data0 (in_0[3]), .sel1 (ctl[3]), .data1
       (in_1[3]), .sel2 (ctl[2]), .data2 (in_2[3]), .sel3 (ctl[1]),
       .data3 (in_3[3]), .sel4 (ctl[0]), .data4 (in_4[3]), .z (z[3]));
  CDN_mux5 g17(.sel0 (ctl[4]), .data0 (in_0[2]), .sel1 (ctl[3]), .data1
       (in_1[2]), .sel2 (ctl[2]), .data2 (in_2[2]), .sel3 (ctl[1]),
       .data3 (in_3[2]), .sel4 (ctl[0]), .data4 (in_4[2]), .z (z[2]));
  CDN_mux5 g18(.sel0 (ctl[4]), .data0 (in_0[1]), .sel1 (ctl[3]), .data1
       (in_1[1]), .sel2 (ctl[2]), .data2 (in_2[1]), .sel3 (ctl[1]),
       .data3 (in_3[1]), .sel4 (ctl[0]), .data4 (in_4[1]), .z (z[1]));
  CDN_mux5 g19(.sel0 (ctl[4]), .data0 (in_0[0]), .sel1 (ctl[3]), .data1
       (in_1[0]), .sel2 (ctl[2]), .data2 (in_2[0]), .sel3 (ctl[1]),
       .data3 (in_3[0]), .sel4 (ctl[0]), .data4 (in_4[0]), .z (z[0]));
endmodule

module fx68k_bmux_299(ctl, in_0, in_1, z);
  input ctl;
  input [9:0] in_0, in_1;
  output [9:0] z;
  wire ctl;
  wire [9:0] in_0, in_1;
  wire [9:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[9]), .data1 (in_1[9]), .z
       (z[9]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[8]), .data1 (in_1[8]), .z
       (z[8]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[7]), .data1 (in_1[7]), .z
       (z[7]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[6]), .data1 (in_1[6]), .z
       (z[6]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g7(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g8(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g9(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g10(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_case_box_83(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_304(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, z);
  input [10:0] ctl;
  input [16:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  output [16:0] z;
  wire [10:0] ctl;
  wire [16:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  wire [16:0] z;
  CDN_mux11 g1(.sel0 (ctl[10]), .data0 (in_0[16]), .sel1 (ctl[9]),
       .data1 (in_1[16]), .sel2 (ctl[8]), .data2 (in_2[16]), .sel3
       (ctl[7]), .data3 (in_3[16]), .sel4 (ctl[6]), .data4 (in_4[16]),
       .sel5 (ctl[5]), .data5 (in_5[16]), .sel6 (ctl[4]), .data6
       (in_6[16]), .sel7 (ctl[3]), .data7 (in_7[16]), .sel8 (ctl[2]),
       .data8 (in_8[16]), .sel9 (ctl[1]), .data9 (in_9[16]), .sel10
       (ctl[0]), .data10 (in_10[16]), .z (z[16]));
  CDN_mux11 g18(.sel0 (ctl[10]), .data0 (in_0[15]), .sel1 (ctl[9]),
       .data1 (in_1[15]), .sel2 (ctl[8]), .data2 (in_2[15]), .sel3
       (ctl[7]), .data3 (in_3[15]), .sel4 (ctl[6]), .data4 (in_4[15]),
       .sel5 (ctl[5]), .data5 (in_5[15]), .sel6 (ctl[4]), .data6
       (in_6[15]), .sel7 (ctl[3]), .data7 (in_7[15]), .sel8 (ctl[2]),
       .data8 (in_8[15]), .sel9 (ctl[1]), .data9 (in_9[15]), .sel10
       (ctl[0]), .data10 (in_10[15]), .z (z[15]));
  CDN_mux11 g19(.sel0 (ctl[10]), .data0 (in_0[14]), .sel1 (ctl[9]),
       .data1 (in_1[14]), .sel2 (ctl[8]), .data2 (in_2[14]), .sel3
       (ctl[7]), .data3 (in_3[14]), .sel4 (ctl[6]), .data4 (in_4[14]),
       .sel5 (ctl[5]), .data5 (in_5[14]), .sel6 (ctl[4]), .data6
       (in_6[14]), .sel7 (ctl[3]), .data7 (in_7[14]), .sel8 (ctl[2]),
       .data8 (in_8[14]), .sel9 (ctl[1]), .data9 (in_9[14]), .sel10
       (ctl[0]), .data10 (in_10[14]), .z (z[14]));
  CDN_mux11 g20(.sel0 (ctl[10]), .data0 (in_0[13]), .sel1 (ctl[9]),
       .data1 (in_1[13]), .sel2 (ctl[8]), .data2 (in_2[13]), .sel3
       (ctl[7]), .data3 (in_3[13]), .sel4 (ctl[6]), .data4 (in_4[13]),
       .sel5 (ctl[5]), .data5 (in_5[13]), .sel6 (ctl[4]), .data6
       (in_6[13]), .sel7 (ctl[3]), .data7 (in_7[13]), .sel8 (ctl[2]),
       .data8 (in_8[13]), .sel9 (ctl[1]), .data9 (in_9[13]), .sel10
       (ctl[0]), .data10 (in_10[13]), .z (z[13]));
  CDN_mux11 g21(.sel0 (ctl[10]), .data0 (in_0[12]), .sel1 (ctl[9]),
       .data1 (in_1[12]), .sel2 (ctl[8]), .data2 (in_2[12]), .sel3
       (ctl[7]), .data3 (in_3[12]), .sel4 (ctl[6]), .data4 (in_4[12]),
       .sel5 (ctl[5]), .data5 (in_5[12]), .sel6 (ctl[4]), .data6
       (in_6[12]), .sel7 (ctl[3]), .data7 (in_7[12]), .sel8 (ctl[2]),
       .data8 (in_8[12]), .sel9 (ctl[1]), .data9 (in_9[12]), .sel10
       (ctl[0]), .data10 (in_10[12]), .z (z[12]));
  CDN_mux11 g22(.sel0 (ctl[10]), .data0 (in_0[11]), .sel1 (ctl[9]),
       .data1 (in_1[11]), .sel2 (ctl[8]), .data2 (in_2[11]), .sel3
       (ctl[7]), .data3 (in_3[11]), .sel4 (ctl[6]), .data4 (in_4[11]),
       .sel5 (ctl[5]), .data5 (in_5[11]), .sel6 (ctl[4]), .data6
       (in_6[11]), .sel7 (ctl[3]), .data7 (in_7[11]), .sel8 (ctl[2]),
       .data8 (in_8[11]), .sel9 (ctl[1]), .data9 (in_9[11]), .sel10
       (ctl[0]), .data10 (in_10[11]), .z (z[11]));
  CDN_mux11 g23(.sel0 (ctl[10]), .data0 (in_0[10]), .sel1 (ctl[9]),
       .data1 (in_1[10]), .sel2 (ctl[8]), .data2 (in_2[10]), .sel3
       (ctl[7]), .data3 (in_3[10]), .sel4 (ctl[6]), .data4 (in_4[10]),
       .sel5 (ctl[5]), .data5 (in_5[10]), .sel6 (ctl[4]), .data6
       (in_6[10]), .sel7 (ctl[3]), .data7 (in_7[10]), .sel8 (ctl[2]),
       .data8 (in_8[10]), .sel9 (ctl[1]), .data9 (in_9[10]), .sel10
       (ctl[0]), .data10 (in_10[10]), .z (z[10]));
  CDN_mux11 g24(.sel0 (ctl[10]), .data0 (in_0[9]), .sel1 (ctl[9]),
       .data1 (in_1[9]), .sel2 (ctl[8]), .data2 (in_2[9]), .sel3
       (ctl[7]), .data3 (in_3[9]), .sel4 (ctl[6]), .data4 (in_4[9]),
       .sel5 (ctl[5]), .data5 (in_5[9]), .sel6 (ctl[4]), .data6
       (in_6[9]), .sel7 (ctl[3]), .data7 (in_7[9]), .sel8 (ctl[2]),
       .data8 (in_8[9]), .sel9 (ctl[1]), .data9 (in_9[9]), .sel10
       (ctl[0]), .data10 (in_10[9]), .z (z[9]));
  CDN_mux11 g25(.sel0 (ctl[10]), .data0 (in_0[8]), .sel1 (ctl[9]),
       .data1 (in_1[8]), .sel2 (ctl[8]), .data2 (in_2[8]), .sel3
       (ctl[7]), .data3 (in_3[8]), .sel4 (ctl[6]), .data4 (in_4[8]),
       .sel5 (ctl[5]), .data5 (in_5[8]), .sel6 (ctl[4]), .data6
       (in_6[8]), .sel7 (ctl[3]), .data7 (in_7[8]), .sel8 (ctl[2]),
       .data8 (in_8[8]), .sel9 (ctl[1]), .data9 (in_9[8]), .sel10
       (ctl[0]), .data10 (in_10[8]), .z (z[8]));
  CDN_mux11 g26(.sel0 (ctl[10]), .data0 (in_0[7]), .sel1 (ctl[9]),
       .data1 (in_1[7]), .sel2 (ctl[8]), .data2 (in_2[7]), .sel3
       (ctl[7]), .data3 (in_3[7]), .sel4 (ctl[6]), .data4 (in_4[7]),
       .sel5 (ctl[5]), .data5 (in_5[7]), .sel6 (ctl[4]), .data6
       (in_6[7]), .sel7 (ctl[3]), .data7 (in_7[7]), .sel8 (ctl[2]),
       .data8 (in_8[7]), .sel9 (ctl[1]), .data9 (in_9[7]), .sel10
       (ctl[0]), .data10 (in_10[7]), .z (z[7]));
  CDN_mux11 g27(.sel0 (ctl[10]), .data0 (in_0[6]), .sel1 (ctl[9]),
       .data1 (in_1[6]), .sel2 (ctl[8]), .data2 (in_2[6]), .sel3
       (ctl[7]), .data3 (in_3[6]), .sel4 (ctl[6]), .data4 (in_4[6]),
       .sel5 (ctl[5]), .data5 (in_5[6]), .sel6 (ctl[4]), .data6
       (in_6[6]), .sel7 (ctl[3]), .data7 (in_7[6]), .sel8 (ctl[2]),
       .data8 (in_8[6]), .sel9 (ctl[1]), .data9 (in_9[6]), .sel10
       (ctl[0]), .data10 (in_10[6]), .z (z[6]));
  CDN_mux11 g28(.sel0 (ctl[10]), .data0 (in_0[5]), .sel1 (ctl[9]),
       .data1 (in_1[5]), .sel2 (ctl[8]), .data2 (in_2[5]), .sel3
       (ctl[7]), .data3 (in_3[5]), .sel4 (ctl[6]), .data4 (in_4[5]),
       .sel5 (ctl[5]), .data5 (in_5[5]), .sel6 (ctl[4]), .data6
       (in_6[5]), .sel7 (ctl[3]), .data7 (in_7[5]), .sel8 (ctl[2]),
       .data8 (in_8[5]), .sel9 (ctl[1]), .data9 (in_9[5]), .sel10
       (ctl[0]), .data10 (in_10[5]), .z (z[5]));
  CDN_mux11 g29(.sel0 (ctl[10]), .data0 (in_0[4]), .sel1 (ctl[9]),
       .data1 (in_1[4]), .sel2 (ctl[8]), .data2 (in_2[4]), .sel3
       (ctl[7]), .data3 (in_3[4]), .sel4 (ctl[6]), .data4 (in_4[4]),
       .sel5 (ctl[5]), .data5 (in_5[4]), .sel6 (ctl[4]), .data6
       (in_6[4]), .sel7 (ctl[3]), .data7 (in_7[4]), .sel8 (ctl[2]),
       .data8 (in_8[4]), .sel9 (ctl[1]), .data9 (in_9[4]), .sel10
       (ctl[0]), .data10 (in_10[4]), .z (z[4]));
  CDN_mux11 g30(.sel0 (ctl[10]), .data0 (in_0[3]), .sel1 (ctl[9]),
       .data1 (in_1[3]), .sel2 (ctl[8]), .data2 (in_2[3]), .sel3
       (ctl[7]), .data3 (in_3[3]), .sel4 (ctl[6]), .data4 (in_4[3]),
       .sel5 (ctl[5]), .data5 (in_5[3]), .sel6 (ctl[4]), .data6
       (in_6[3]), .sel7 (ctl[3]), .data7 (in_7[3]), .sel8 (ctl[2]),
       .data8 (in_8[3]), .sel9 (ctl[1]), .data9 (in_9[3]), .sel10
       (ctl[0]), .data10 (in_10[3]), .z (z[3]));
  CDN_mux11 g31(.sel0 (ctl[10]), .data0 (in_0[2]), .sel1 (ctl[9]),
       .data1 (in_1[2]), .sel2 (ctl[8]), .data2 (in_2[2]), .sel3
       (ctl[7]), .data3 (in_3[2]), .sel4 (ctl[6]), .data4 (in_4[2]),
       .sel5 (ctl[5]), .data5 (in_5[2]), .sel6 (ctl[4]), .data6
       (in_6[2]), .sel7 (ctl[3]), .data7 (in_7[2]), .sel8 (ctl[2]),
       .data8 (in_8[2]), .sel9 (ctl[1]), .data9 (in_9[2]), .sel10
       (ctl[0]), .data10 (in_10[2]), .z (z[2]));
  CDN_mux11 g32(.sel0 (ctl[10]), .data0 (in_0[1]), .sel1 (ctl[9]),
       .data1 (in_1[1]), .sel2 (ctl[8]), .data2 (in_2[1]), .sel3
       (ctl[7]), .data3 (in_3[1]), .sel4 (ctl[6]), .data4 (in_4[1]),
       .sel5 (ctl[5]), .data5 (in_5[1]), .sel6 (ctl[4]), .data6
       (in_6[1]), .sel7 (ctl[3]), .data7 (in_7[1]), .sel8 (ctl[2]),
       .data8 (in_8[1]), .sel9 (ctl[1]), .data9 (in_9[1]), .sel10
       (ctl[0]), .data10 (in_10[1]), .z (z[1]));
  CDN_mux11 g33(.sel0 (ctl[10]), .data0 (in_0[0]), .sel1 (ctl[9]),
       .data1 (in_1[0]), .sel2 (ctl[8]), .data2 (in_2[0]), .sel3
       (ctl[7]), .data3 (in_3[0]), .sel4 (ctl[6]), .data4 (in_4[0]),
       .sel5 (ctl[5]), .data5 (in_5[0]), .sel6 (ctl[4]), .data6
       (in_6[0]), .sel7 (ctl[3]), .data7 (in_7[0]), .sel8 (ctl[2]),
       .data8 (in_8[0]), .sel9 (ctl[1]), .data9 (in_9[0]), .sel10
       (ctl[0]), .data10 (in_10[0]), .z (z[0]));
endmodule

module fx68k_case_box_86(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_320(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, z);
  input [10:0] ctl;
  input [13:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  output [13:0] z;
  wire [10:0] ctl;
  wire [13:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  wire [13:0] z;
  CDN_mux11 g1(.sel0 (ctl[10]), .data0 (in_0[13]), .sel1 (ctl[9]),
       .data1 (in_1[13]), .sel2 (ctl[8]), .data2 (in_2[13]), .sel3
       (ctl[7]), .data3 (in_3[13]), .sel4 (ctl[6]), .data4 (in_4[13]),
       .sel5 (ctl[5]), .data5 (in_5[13]), .sel6 (ctl[4]), .data6
       (in_6[13]), .sel7 (ctl[3]), .data7 (in_7[13]), .sel8 (ctl[2]),
       .data8 (in_8[13]), .sel9 (ctl[1]), .data9 (in_9[13]), .sel10
       (ctl[0]), .data10 (in_10[13]), .z (z[13]));
  CDN_mux11 g15(.sel0 (ctl[10]), .data0 (in_0[12]), .sel1 (ctl[9]),
       .data1 (in_1[12]), .sel2 (ctl[8]), .data2 (in_2[12]), .sel3
       (ctl[7]), .data3 (in_3[12]), .sel4 (ctl[6]), .data4 (in_4[12]),
       .sel5 (ctl[5]), .data5 (in_5[12]), .sel6 (ctl[4]), .data6
       (in_6[12]), .sel7 (ctl[3]), .data7 (in_7[12]), .sel8 (ctl[2]),
       .data8 (in_8[12]), .sel9 (ctl[1]), .data9 (in_9[12]), .sel10
       (ctl[0]), .data10 (in_10[12]), .z (z[12]));
  CDN_mux11 g16(.sel0 (ctl[10]), .data0 (in_0[11]), .sel1 (ctl[9]),
       .data1 (in_1[11]), .sel2 (ctl[8]), .data2 (in_2[11]), .sel3
       (ctl[7]), .data3 (in_3[11]), .sel4 (ctl[6]), .data4 (in_4[11]),
       .sel5 (ctl[5]), .data5 (in_5[11]), .sel6 (ctl[4]), .data6
       (in_6[11]), .sel7 (ctl[3]), .data7 (in_7[11]), .sel8 (ctl[2]),
       .data8 (in_8[11]), .sel9 (ctl[1]), .data9 (in_9[11]), .sel10
       (ctl[0]), .data10 (in_10[11]), .z (z[11]));
  CDN_mux11 g17(.sel0 (ctl[10]), .data0 (in_0[10]), .sel1 (ctl[9]),
       .data1 (in_1[10]), .sel2 (ctl[8]), .data2 (in_2[10]), .sel3
       (ctl[7]), .data3 (in_3[10]), .sel4 (ctl[6]), .data4 (in_4[10]),
       .sel5 (ctl[5]), .data5 (in_5[10]), .sel6 (ctl[4]), .data6
       (in_6[10]), .sel7 (ctl[3]), .data7 (in_7[10]), .sel8 (ctl[2]),
       .data8 (in_8[10]), .sel9 (ctl[1]), .data9 (in_9[10]), .sel10
       (ctl[0]), .data10 (in_10[10]), .z (z[10]));
  CDN_mux11 g18(.sel0 (ctl[10]), .data0 (in_0[9]), .sel1 (ctl[9]),
       .data1 (in_1[9]), .sel2 (ctl[8]), .data2 (in_2[9]), .sel3
       (ctl[7]), .data3 (in_3[9]), .sel4 (ctl[6]), .data4 (in_4[9]),
       .sel5 (ctl[5]), .data5 (in_5[9]), .sel6 (ctl[4]), .data6
       (in_6[9]), .sel7 (ctl[3]), .data7 (in_7[9]), .sel8 (ctl[2]),
       .data8 (in_8[9]), .sel9 (ctl[1]), .data9 (in_9[9]), .sel10
       (ctl[0]), .data10 (in_10[9]), .z (z[9]));
  CDN_mux11 g19(.sel0 (ctl[10]), .data0 (in_0[8]), .sel1 (ctl[9]),
       .data1 (in_1[8]), .sel2 (ctl[8]), .data2 (in_2[8]), .sel3
       (ctl[7]), .data3 (in_3[8]), .sel4 (ctl[6]), .data4 (in_4[8]),
       .sel5 (ctl[5]), .data5 (in_5[8]), .sel6 (ctl[4]), .data6
       (in_6[8]), .sel7 (ctl[3]), .data7 (in_7[8]), .sel8 (ctl[2]),
       .data8 (in_8[8]), .sel9 (ctl[1]), .data9 (in_9[8]), .sel10
       (ctl[0]), .data10 (in_10[8]), .z (z[8]));
  CDN_mux11 g20(.sel0 (ctl[10]), .data0 (in_0[7]), .sel1 (ctl[9]),
       .data1 (in_1[7]), .sel2 (ctl[8]), .data2 (in_2[7]), .sel3
       (ctl[7]), .data3 (in_3[7]), .sel4 (ctl[6]), .data4 (in_4[7]),
       .sel5 (ctl[5]), .data5 (in_5[7]), .sel6 (ctl[4]), .data6
       (in_6[7]), .sel7 (ctl[3]), .data7 (in_7[7]), .sel8 (ctl[2]),
       .data8 (in_8[7]), .sel9 (ctl[1]), .data9 (in_9[7]), .sel10
       (ctl[0]), .data10 (in_10[7]), .z (z[7]));
  CDN_mux11 g21(.sel0 (ctl[10]), .data0 (in_0[6]), .sel1 (ctl[9]),
       .data1 (in_1[6]), .sel2 (ctl[8]), .data2 (in_2[6]), .sel3
       (ctl[7]), .data3 (in_3[6]), .sel4 (ctl[6]), .data4 (in_4[6]),
       .sel5 (ctl[5]), .data5 (in_5[6]), .sel6 (ctl[4]), .data6
       (in_6[6]), .sel7 (ctl[3]), .data7 (in_7[6]), .sel8 (ctl[2]),
       .data8 (in_8[6]), .sel9 (ctl[1]), .data9 (in_9[6]), .sel10
       (ctl[0]), .data10 (in_10[6]), .z (z[6]));
  CDN_mux11 g22(.sel0 (ctl[10]), .data0 (in_0[5]), .sel1 (ctl[9]),
       .data1 (in_1[5]), .sel2 (ctl[8]), .data2 (in_2[5]), .sel3
       (ctl[7]), .data3 (in_3[5]), .sel4 (ctl[6]), .data4 (in_4[5]),
       .sel5 (ctl[5]), .data5 (in_5[5]), .sel6 (ctl[4]), .data6
       (in_6[5]), .sel7 (ctl[3]), .data7 (in_7[5]), .sel8 (ctl[2]),
       .data8 (in_8[5]), .sel9 (ctl[1]), .data9 (in_9[5]), .sel10
       (ctl[0]), .data10 (in_10[5]), .z (z[5]));
  CDN_mux11 g23(.sel0 (ctl[10]), .data0 (in_0[4]), .sel1 (ctl[9]),
       .data1 (in_1[4]), .sel2 (ctl[8]), .data2 (in_2[4]), .sel3
       (ctl[7]), .data3 (in_3[4]), .sel4 (ctl[6]), .data4 (in_4[4]),
       .sel5 (ctl[5]), .data5 (in_5[4]), .sel6 (ctl[4]), .data6
       (in_6[4]), .sel7 (ctl[3]), .data7 (in_7[4]), .sel8 (ctl[2]),
       .data8 (in_8[4]), .sel9 (ctl[1]), .data9 (in_9[4]), .sel10
       (ctl[0]), .data10 (in_10[4]), .z (z[4]));
  CDN_mux11 g24(.sel0 (ctl[10]), .data0 (in_0[3]), .sel1 (ctl[9]),
       .data1 (in_1[3]), .sel2 (ctl[8]), .data2 (in_2[3]), .sel3
       (ctl[7]), .data3 (in_3[3]), .sel4 (ctl[6]), .data4 (in_4[3]),
       .sel5 (ctl[5]), .data5 (in_5[3]), .sel6 (ctl[4]), .data6
       (in_6[3]), .sel7 (ctl[3]), .data7 (in_7[3]), .sel8 (ctl[2]),
       .data8 (in_8[3]), .sel9 (ctl[1]), .data9 (in_9[3]), .sel10
       (ctl[0]), .data10 (in_10[3]), .z (z[3]));
  CDN_mux11 g25(.sel0 (ctl[10]), .data0 (in_0[2]), .sel1 (ctl[9]),
       .data1 (in_1[2]), .sel2 (ctl[8]), .data2 (in_2[2]), .sel3
       (ctl[7]), .data3 (in_3[2]), .sel4 (ctl[6]), .data4 (in_4[2]),
       .sel5 (ctl[5]), .data5 (in_5[2]), .sel6 (ctl[4]), .data6
       (in_6[2]), .sel7 (ctl[3]), .data7 (in_7[2]), .sel8 (ctl[2]),
       .data8 (in_8[2]), .sel9 (ctl[1]), .data9 (in_9[2]), .sel10
       (ctl[0]), .data10 (in_10[2]), .z (z[2]));
  CDN_mux11 g26(.sel0 (ctl[10]), .data0 (in_0[1]), .sel1 (ctl[9]),
       .data1 (in_1[1]), .sel2 (ctl[8]), .data2 (in_2[1]), .sel3
       (ctl[7]), .data3 (in_3[1]), .sel4 (ctl[6]), .data4 (in_4[1]),
       .sel5 (ctl[5]), .data5 (in_5[1]), .sel6 (ctl[4]), .data6
       (in_6[1]), .sel7 (ctl[3]), .data7 (in_7[1]), .sel8 (ctl[2]),
       .data8 (in_8[1]), .sel9 (ctl[1]), .data9 (in_9[1]), .sel10
       (ctl[0]), .data10 (in_10[1]), .z (z[1]));
  CDN_mux11 g27(.sel0 (ctl[10]), .data0 (in_0[0]), .sel1 (ctl[9]),
       .data1 (in_1[0]), .sel2 (ctl[8]), .data2 (in_2[0]), .sel3
       (ctl[7]), .data3 (in_3[0]), .sel4 (ctl[6]), .data4 (in_4[0]),
       .sel5 (ctl[5]), .data5 (in_5[0]), .sel6 (ctl[4]), .data6
       (in_6[0]), .sel7 (ctl[3]), .data7 (in_7[0]), .sel8 (ctl[2]),
       .data8 (in_8[0]), .sel9 (ctl[1]), .data9 (in_9[0]), .sel10
       (ctl[0]), .data10 (in_10[0]), .z (z[0]));
endmodule

module fx68k_case_box_89(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_92(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_346(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, z);
  input [10:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  output [15:0] z;
  wire [10:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  wire [15:0] z;
  CDN_mux11 g1(.sel0 (ctl[10]), .data0 (in_0[15]), .sel1 (ctl[9]),
       .data1 (in_1[15]), .sel2 (ctl[8]), .data2 (in_2[15]), .sel3
       (ctl[7]), .data3 (in_3[15]), .sel4 (ctl[6]), .data4 (in_4[15]),
       .sel5 (ctl[5]), .data5 (in_5[15]), .sel6 (ctl[4]), .data6
       (in_6[15]), .sel7 (ctl[3]), .data7 (in_7[15]), .sel8 (ctl[2]),
       .data8 (in_8[15]), .sel9 (ctl[1]), .data9 (in_9[15]), .sel10
       (ctl[0]), .data10 (in_10[15]), .z (z[15]));
  CDN_mux11 g17(.sel0 (ctl[10]), .data0 (in_0[14]), .sel1 (ctl[9]),
       .data1 (in_1[14]), .sel2 (ctl[8]), .data2 (in_2[14]), .sel3
       (ctl[7]), .data3 (in_3[14]), .sel4 (ctl[6]), .data4 (in_4[14]),
       .sel5 (ctl[5]), .data5 (in_5[14]), .sel6 (ctl[4]), .data6
       (in_6[14]), .sel7 (ctl[3]), .data7 (in_7[14]), .sel8 (ctl[2]),
       .data8 (in_8[14]), .sel9 (ctl[1]), .data9 (in_9[14]), .sel10
       (ctl[0]), .data10 (in_10[14]), .z (z[14]));
  CDN_mux11 g18(.sel0 (ctl[10]), .data0 (in_0[13]), .sel1 (ctl[9]),
       .data1 (in_1[13]), .sel2 (ctl[8]), .data2 (in_2[13]), .sel3
       (ctl[7]), .data3 (in_3[13]), .sel4 (ctl[6]), .data4 (in_4[13]),
       .sel5 (ctl[5]), .data5 (in_5[13]), .sel6 (ctl[4]), .data6
       (in_6[13]), .sel7 (ctl[3]), .data7 (in_7[13]), .sel8 (ctl[2]),
       .data8 (in_8[13]), .sel9 (ctl[1]), .data9 (in_9[13]), .sel10
       (ctl[0]), .data10 (in_10[13]), .z (z[13]));
  CDN_mux11 g19(.sel0 (ctl[10]), .data0 (in_0[12]), .sel1 (ctl[9]),
       .data1 (in_1[12]), .sel2 (ctl[8]), .data2 (in_2[12]), .sel3
       (ctl[7]), .data3 (in_3[12]), .sel4 (ctl[6]), .data4 (in_4[12]),
       .sel5 (ctl[5]), .data5 (in_5[12]), .sel6 (ctl[4]), .data6
       (in_6[12]), .sel7 (ctl[3]), .data7 (in_7[12]), .sel8 (ctl[2]),
       .data8 (in_8[12]), .sel9 (ctl[1]), .data9 (in_9[12]), .sel10
       (ctl[0]), .data10 (in_10[12]), .z (z[12]));
  CDN_mux11 g20(.sel0 (ctl[10]), .data0 (in_0[11]), .sel1 (ctl[9]),
       .data1 (in_1[11]), .sel2 (ctl[8]), .data2 (in_2[11]), .sel3
       (ctl[7]), .data3 (in_3[11]), .sel4 (ctl[6]), .data4 (in_4[11]),
       .sel5 (ctl[5]), .data5 (in_5[11]), .sel6 (ctl[4]), .data6
       (in_6[11]), .sel7 (ctl[3]), .data7 (in_7[11]), .sel8 (ctl[2]),
       .data8 (in_8[11]), .sel9 (ctl[1]), .data9 (in_9[11]), .sel10
       (ctl[0]), .data10 (in_10[11]), .z (z[11]));
  CDN_mux11 g21(.sel0 (ctl[10]), .data0 (in_0[10]), .sel1 (ctl[9]),
       .data1 (in_1[10]), .sel2 (ctl[8]), .data2 (in_2[10]), .sel3
       (ctl[7]), .data3 (in_3[10]), .sel4 (ctl[6]), .data4 (in_4[10]),
       .sel5 (ctl[5]), .data5 (in_5[10]), .sel6 (ctl[4]), .data6
       (in_6[10]), .sel7 (ctl[3]), .data7 (in_7[10]), .sel8 (ctl[2]),
       .data8 (in_8[10]), .sel9 (ctl[1]), .data9 (in_9[10]), .sel10
       (ctl[0]), .data10 (in_10[10]), .z (z[10]));
  CDN_mux11 g22(.sel0 (ctl[10]), .data0 (in_0[9]), .sel1 (ctl[9]),
       .data1 (in_1[9]), .sel2 (ctl[8]), .data2 (in_2[9]), .sel3
       (ctl[7]), .data3 (in_3[9]), .sel4 (ctl[6]), .data4 (in_4[9]),
       .sel5 (ctl[5]), .data5 (in_5[9]), .sel6 (ctl[4]), .data6
       (in_6[9]), .sel7 (ctl[3]), .data7 (in_7[9]), .sel8 (ctl[2]),
       .data8 (in_8[9]), .sel9 (ctl[1]), .data9 (in_9[9]), .sel10
       (ctl[0]), .data10 (in_10[9]), .z (z[9]));
  CDN_mux11 g23(.sel0 (ctl[10]), .data0 (in_0[8]), .sel1 (ctl[9]),
       .data1 (in_1[8]), .sel2 (ctl[8]), .data2 (in_2[8]), .sel3
       (ctl[7]), .data3 (in_3[8]), .sel4 (ctl[6]), .data4 (in_4[8]),
       .sel5 (ctl[5]), .data5 (in_5[8]), .sel6 (ctl[4]), .data6
       (in_6[8]), .sel7 (ctl[3]), .data7 (in_7[8]), .sel8 (ctl[2]),
       .data8 (in_8[8]), .sel9 (ctl[1]), .data9 (in_9[8]), .sel10
       (ctl[0]), .data10 (in_10[8]), .z (z[8]));
  CDN_mux11 g24(.sel0 (ctl[10]), .data0 (in_0[7]), .sel1 (ctl[9]),
       .data1 (in_1[7]), .sel2 (ctl[8]), .data2 (in_2[7]), .sel3
       (ctl[7]), .data3 (in_3[7]), .sel4 (ctl[6]), .data4 (in_4[7]),
       .sel5 (ctl[5]), .data5 (in_5[7]), .sel6 (ctl[4]), .data6
       (in_6[7]), .sel7 (ctl[3]), .data7 (in_7[7]), .sel8 (ctl[2]),
       .data8 (in_8[7]), .sel9 (ctl[1]), .data9 (in_9[7]), .sel10
       (ctl[0]), .data10 (in_10[7]), .z (z[7]));
  CDN_mux11 g25(.sel0 (ctl[10]), .data0 (in_0[6]), .sel1 (ctl[9]),
       .data1 (in_1[6]), .sel2 (ctl[8]), .data2 (in_2[6]), .sel3
       (ctl[7]), .data3 (in_3[6]), .sel4 (ctl[6]), .data4 (in_4[6]),
       .sel5 (ctl[5]), .data5 (in_5[6]), .sel6 (ctl[4]), .data6
       (in_6[6]), .sel7 (ctl[3]), .data7 (in_7[6]), .sel8 (ctl[2]),
       .data8 (in_8[6]), .sel9 (ctl[1]), .data9 (in_9[6]), .sel10
       (ctl[0]), .data10 (in_10[6]), .z (z[6]));
  CDN_mux11 g26(.sel0 (ctl[10]), .data0 (in_0[5]), .sel1 (ctl[9]),
       .data1 (in_1[5]), .sel2 (ctl[8]), .data2 (in_2[5]), .sel3
       (ctl[7]), .data3 (in_3[5]), .sel4 (ctl[6]), .data4 (in_4[5]),
       .sel5 (ctl[5]), .data5 (in_5[5]), .sel6 (ctl[4]), .data6
       (in_6[5]), .sel7 (ctl[3]), .data7 (in_7[5]), .sel8 (ctl[2]),
       .data8 (in_8[5]), .sel9 (ctl[1]), .data9 (in_9[5]), .sel10
       (ctl[0]), .data10 (in_10[5]), .z (z[5]));
  CDN_mux11 g27(.sel0 (ctl[10]), .data0 (in_0[4]), .sel1 (ctl[9]),
       .data1 (in_1[4]), .sel2 (ctl[8]), .data2 (in_2[4]), .sel3
       (ctl[7]), .data3 (in_3[4]), .sel4 (ctl[6]), .data4 (in_4[4]),
       .sel5 (ctl[5]), .data5 (in_5[4]), .sel6 (ctl[4]), .data6
       (in_6[4]), .sel7 (ctl[3]), .data7 (in_7[4]), .sel8 (ctl[2]),
       .data8 (in_8[4]), .sel9 (ctl[1]), .data9 (in_9[4]), .sel10
       (ctl[0]), .data10 (in_10[4]), .z (z[4]));
  CDN_mux11 g28(.sel0 (ctl[10]), .data0 (in_0[3]), .sel1 (ctl[9]),
       .data1 (in_1[3]), .sel2 (ctl[8]), .data2 (in_2[3]), .sel3
       (ctl[7]), .data3 (in_3[3]), .sel4 (ctl[6]), .data4 (in_4[3]),
       .sel5 (ctl[5]), .data5 (in_5[3]), .sel6 (ctl[4]), .data6
       (in_6[3]), .sel7 (ctl[3]), .data7 (in_7[3]), .sel8 (ctl[2]),
       .data8 (in_8[3]), .sel9 (ctl[1]), .data9 (in_9[3]), .sel10
       (ctl[0]), .data10 (in_10[3]), .z (z[3]));
  CDN_mux11 g29(.sel0 (ctl[10]), .data0 (in_0[2]), .sel1 (ctl[9]),
       .data1 (in_1[2]), .sel2 (ctl[8]), .data2 (in_2[2]), .sel3
       (ctl[7]), .data3 (in_3[2]), .sel4 (ctl[6]), .data4 (in_4[2]),
       .sel5 (ctl[5]), .data5 (in_5[2]), .sel6 (ctl[4]), .data6
       (in_6[2]), .sel7 (ctl[3]), .data7 (in_7[2]), .sel8 (ctl[2]),
       .data8 (in_8[2]), .sel9 (ctl[1]), .data9 (in_9[2]), .sel10
       (ctl[0]), .data10 (in_10[2]), .z (z[2]));
  CDN_mux11 g30(.sel0 (ctl[10]), .data0 (in_0[1]), .sel1 (ctl[9]),
       .data1 (in_1[1]), .sel2 (ctl[8]), .data2 (in_2[1]), .sel3
       (ctl[7]), .data3 (in_3[1]), .sel4 (ctl[6]), .data4 (in_4[1]),
       .sel5 (ctl[5]), .data5 (in_5[1]), .sel6 (ctl[4]), .data6
       (in_6[1]), .sel7 (ctl[3]), .data7 (in_7[1]), .sel8 (ctl[2]),
       .data8 (in_8[1]), .sel9 (ctl[1]), .data9 (in_9[1]), .sel10
       (ctl[0]), .data10 (in_10[1]), .z (z[1]));
  CDN_mux11 g31(.sel0 (ctl[10]), .data0 (in_0[0]), .sel1 (ctl[9]),
       .data1 (in_1[0]), .sel2 (ctl[8]), .data2 (in_2[0]), .sel3
       (ctl[7]), .data3 (in_3[0]), .sel4 (ctl[6]), .data4 (in_4[0]),
       .sel5 (ctl[5]), .data5 (in_5[0]), .sel6 (ctl[4]), .data6
       (in_6[0]), .sel7 (ctl[3]), .data7 (in_7[0]), .sel8 (ctl[2]),
       .data8 (in_8[0]), .sel9 (ctl[1]), .data9 (in_9[0]), .sel10
       (ctl[0]), .data10 (in_10[0]), .z (z[0]));
endmodule

module fx68k_case_box_95(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_361(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, z);
  input [10:0] ctl;
  input [12:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  output [12:0] z;
  wire [10:0] ctl;
  wire [12:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  wire [12:0] z;
  CDN_mux11 g1(.sel0 (ctl[10]), .data0 (in_0[12]), .sel1 (ctl[9]),
       .data1 (in_1[12]), .sel2 (ctl[8]), .data2 (in_2[12]), .sel3
       (ctl[7]), .data3 (in_3[12]), .sel4 (ctl[6]), .data4 (in_4[12]),
       .sel5 (ctl[5]), .data5 (in_5[12]), .sel6 (ctl[4]), .data6
       (in_6[12]), .sel7 (ctl[3]), .data7 (in_7[12]), .sel8 (ctl[2]),
       .data8 (in_8[12]), .sel9 (ctl[1]), .data9 (in_9[12]), .sel10
       (ctl[0]), .data10 (in_10[12]), .z (z[12]));
  CDN_mux11 g14(.sel0 (ctl[10]), .data0 (in_0[11]), .sel1 (ctl[9]),
       .data1 (in_1[11]), .sel2 (ctl[8]), .data2 (in_2[11]), .sel3
       (ctl[7]), .data3 (in_3[11]), .sel4 (ctl[6]), .data4 (in_4[11]),
       .sel5 (ctl[5]), .data5 (in_5[11]), .sel6 (ctl[4]), .data6
       (in_6[11]), .sel7 (ctl[3]), .data7 (in_7[11]), .sel8 (ctl[2]),
       .data8 (in_8[11]), .sel9 (ctl[1]), .data9 (in_9[11]), .sel10
       (ctl[0]), .data10 (in_10[11]), .z (z[11]));
  CDN_mux11 g15(.sel0 (ctl[10]), .data0 (in_0[10]), .sel1 (ctl[9]),
       .data1 (in_1[10]), .sel2 (ctl[8]), .data2 (in_2[10]), .sel3
       (ctl[7]), .data3 (in_3[10]), .sel4 (ctl[6]), .data4 (in_4[10]),
       .sel5 (ctl[5]), .data5 (in_5[10]), .sel6 (ctl[4]), .data6
       (in_6[10]), .sel7 (ctl[3]), .data7 (in_7[10]), .sel8 (ctl[2]),
       .data8 (in_8[10]), .sel9 (ctl[1]), .data9 (in_9[10]), .sel10
       (ctl[0]), .data10 (in_10[10]), .z (z[10]));
  CDN_mux11 g16(.sel0 (ctl[10]), .data0 (in_0[9]), .sel1 (ctl[9]),
       .data1 (in_1[9]), .sel2 (ctl[8]), .data2 (in_2[9]), .sel3
       (ctl[7]), .data3 (in_3[9]), .sel4 (ctl[6]), .data4 (in_4[9]),
       .sel5 (ctl[5]), .data5 (in_5[9]), .sel6 (ctl[4]), .data6
       (in_6[9]), .sel7 (ctl[3]), .data7 (in_7[9]), .sel8 (ctl[2]),
       .data8 (in_8[9]), .sel9 (ctl[1]), .data9 (in_9[9]), .sel10
       (ctl[0]), .data10 (in_10[9]), .z (z[9]));
  CDN_mux11 g17(.sel0 (ctl[10]), .data0 (in_0[8]), .sel1 (ctl[9]),
       .data1 (in_1[8]), .sel2 (ctl[8]), .data2 (in_2[8]), .sel3
       (ctl[7]), .data3 (in_3[8]), .sel4 (ctl[6]), .data4 (in_4[8]),
       .sel5 (ctl[5]), .data5 (in_5[8]), .sel6 (ctl[4]), .data6
       (in_6[8]), .sel7 (ctl[3]), .data7 (in_7[8]), .sel8 (ctl[2]),
       .data8 (in_8[8]), .sel9 (ctl[1]), .data9 (in_9[8]), .sel10
       (ctl[0]), .data10 (in_10[8]), .z (z[8]));
  CDN_mux11 g18(.sel0 (ctl[10]), .data0 (in_0[7]), .sel1 (ctl[9]),
       .data1 (in_1[7]), .sel2 (ctl[8]), .data2 (in_2[7]), .sel3
       (ctl[7]), .data3 (in_3[7]), .sel4 (ctl[6]), .data4 (in_4[7]),
       .sel5 (ctl[5]), .data5 (in_5[7]), .sel6 (ctl[4]), .data6
       (in_6[7]), .sel7 (ctl[3]), .data7 (in_7[7]), .sel8 (ctl[2]),
       .data8 (in_8[7]), .sel9 (ctl[1]), .data9 (in_9[7]), .sel10
       (ctl[0]), .data10 (in_10[7]), .z (z[7]));
  CDN_mux11 g19(.sel0 (ctl[10]), .data0 (in_0[6]), .sel1 (ctl[9]),
       .data1 (in_1[6]), .sel2 (ctl[8]), .data2 (in_2[6]), .sel3
       (ctl[7]), .data3 (in_3[6]), .sel4 (ctl[6]), .data4 (in_4[6]),
       .sel5 (ctl[5]), .data5 (in_5[6]), .sel6 (ctl[4]), .data6
       (in_6[6]), .sel7 (ctl[3]), .data7 (in_7[6]), .sel8 (ctl[2]),
       .data8 (in_8[6]), .sel9 (ctl[1]), .data9 (in_9[6]), .sel10
       (ctl[0]), .data10 (in_10[6]), .z (z[6]));
  CDN_mux11 g20(.sel0 (ctl[10]), .data0 (in_0[5]), .sel1 (ctl[9]),
       .data1 (in_1[5]), .sel2 (ctl[8]), .data2 (in_2[5]), .sel3
       (ctl[7]), .data3 (in_3[5]), .sel4 (ctl[6]), .data4 (in_4[5]),
       .sel5 (ctl[5]), .data5 (in_5[5]), .sel6 (ctl[4]), .data6
       (in_6[5]), .sel7 (ctl[3]), .data7 (in_7[5]), .sel8 (ctl[2]),
       .data8 (in_8[5]), .sel9 (ctl[1]), .data9 (in_9[5]), .sel10
       (ctl[0]), .data10 (in_10[5]), .z (z[5]));
  CDN_mux11 g21(.sel0 (ctl[10]), .data0 (in_0[4]), .sel1 (ctl[9]),
       .data1 (in_1[4]), .sel2 (ctl[8]), .data2 (in_2[4]), .sel3
       (ctl[7]), .data3 (in_3[4]), .sel4 (ctl[6]), .data4 (in_4[4]),
       .sel5 (ctl[5]), .data5 (in_5[4]), .sel6 (ctl[4]), .data6
       (in_6[4]), .sel7 (ctl[3]), .data7 (in_7[4]), .sel8 (ctl[2]),
       .data8 (in_8[4]), .sel9 (ctl[1]), .data9 (in_9[4]), .sel10
       (ctl[0]), .data10 (in_10[4]), .z (z[4]));
  CDN_mux11 g22(.sel0 (ctl[10]), .data0 (in_0[3]), .sel1 (ctl[9]),
       .data1 (in_1[3]), .sel2 (ctl[8]), .data2 (in_2[3]), .sel3
       (ctl[7]), .data3 (in_3[3]), .sel4 (ctl[6]), .data4 (in_4[3]),
       .sel5 (ctl[5]), .data5 (in_5[3]), .sel6 (ctl[4]), .data6
       (in_6[3]), .sel7 (ctl[3]), .data7 (in_7[3]), .sel8 (ctl[2]),
       .data8 (in_8[3]), .sel9 (ctl[1]), .data9 (in_9[3]), .sel10
       (ctl[0]), .data10 (in_10[3]), .z (z[3]));
  CDN_mux11 g23(.sel0 (ctl[10]), .data0 (in_0[2]), .sel1 (ctl[9]),
       .data1 (in_1[2]), .sel2 (ctl[8]), .data2 (in_2[2]), .sel3
       (ctl[7]), .data3 (in_3[2]), .sel4 (ctl[6]), .data4 (in_4[2]),
       .sel5 (ctl[5]), .data5 (in_5[2]), .sel6 (ctl[4]), .data6
       (in_6[2]), .sel7 (ctl[3]), .data7 (in_7[2]), .sel8 (ctl[2]),
       .data8 (in_8[2]), .sel9 (ctl[1]), .data9 (in_9[2]), .sel10
       (ctl[0]), .data10 (in_10[2]), .z (z[2]));
  CDN_mux11 g24(.sel0 (ctl[10]), .data0 (in_0[1]), .sel1 (ctl[9]),
       .data1 (in_1[1]), .sel2 (ctl[8]), .data2 (in_2[1]), .sel3
       (ctl[7]), .data3 (in_3[1]), .sel4 (ctl[6]), .data4 (in_4[1]),
       .sel5 (ctl[5]), .data5 (in_5[1]), .sel6 (ctl[4]), .data6
       (in_6[1]), .sel7 (ctl[3]), .data7 (in_7[1]), .sel8 (ctl[2]),
       .data8 (in_8[1]), .sel9 (ctl[1]), .data9 (in_9[1]), .sel10
       (ctl[0]), .data10 (in_10[1]), .z (z[1]));
  CDN_mux11 g25(.sel0 (ctl[10]), .data0 (in_0[0]), .sel1 (ctl[9]),
       .data1 (in_1[0]), .sel2 (ctl[8]), .data2 (in_2[0]), .sel3
       (ctl[7]), .data3 (in_3[0]), .sel4 (ctl[6]), .data4 (in_4[0]),
       .sel5 (ctl[5]), .data5 (in_5[0]), .sel6 (ctl[4]), .data6
       (in_6[0]), .sel7 (ctl[3]), .data7 (in_7[0]), .sel8 (ctl[2]),
       .data8 (in_8[0]), .sel9 (ctl[1]), .data9 (in_9[0]), .sel10
       (ctl[0]), .data10 (in_10[0]), .z (z[0]));
endmodule

module fx68k_case_box_98(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_101(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_104(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_110(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_424(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  output [15:0] z;
  wire [11:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  wire [15:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[15]), .sel1 (ctl[10]),
       .data1 (in_1[15]), .sel2 (ctl[9]), .data2 (in_2[15]), .sel3
       (ctl[8]), .data3 (in_3[15]), .sel4 (ctl[7]), .data4 (in_4[15]),
       .sel5 (ctl[6]), .data5 (in_5[15]), .sel6 (ctl[5]), .data6
       (in_6[15]), .sel7 (ctl[4]), .data7 (in_7[15]), .sel8 (ctl[3]),
       .data8 (in_8[15]), .sel9 (ctl[2]), .data9 (in_9[15]), .sel10
       (ctl[1]), .data10 (in_10[15]), .sel11 (ctl[0]), .data11
       (in_11[15]), .z (z[15]));
  CDN_mux12 g17(.sel0 (ctl[11]), .data0 (in_0[14]), .sel1 (ctl[10]),
       .data1 (in_1[14]), .sel2 (ctl[9]), .data2 (in_2[14]), .sel3
       (ctl[8]), .data3 (in_3[14]), .sel4 (ctl[7]), .data4 (in_4[14]),
       .sel5 (ctl[6]), .data5 (in_5[14]), .sel6 (ctl[5]), .data6
       (in_6[14]), .sel7 (ctl[4]), .data7 (in_7[14]), .sel8 (ctl[3]),
       .data8 (in_8[14]), .sel9 (ctl[2]), .data9 (in_9[14]), .sel10
       (ctl[1]), .data10 (in_10[14]), .sel11 (ctl[0]), .data11
       (in_11[14]), .z (z[14]));
  CDN_mux12 g18(.sel0 (ctl[11]), .data0 (in_0[13]), .sel1 (ctl[10]),
       .data1 (in_1[13]), .sel2 (ctl[9]), .data2 (in_2[13]), .sel3
       (ctl[8]), .data3 (in_3[13]), .sel4 (ctl[7]), .data4 (in_4[13]),
       .sel5 (ctl[6]), .data5 (in_5[13]), .sel6 (ctl[5]), .data6
       (in_6[13]), .sel7 (ctl[4]), .data7 (in_7[13]), .sel8 (ctl[3]),
       .data8 (in_8[13]), .sel9 (ctl[2]), .data9 (in_9[13]), .sel10
       (ctl[1]), .data10 (in_10[13]), .sel11 (ctl[0]), .data11
       (in_11[13]), .z (z[13]));
  CDN_mux12 g19(.sel0 (ctl[11]), .data0 (in_0[12]), .sel1 (ctl[10]),
       .data1 (in_1[12]), .sel2 (ctl[9]), .data2 (in_2[12]), .sel3
       (ctl[8]), .data3 (in_3[12]), .sel4 (ctl[7]), .data4 (in_4[12]),
       .sel5 (ctl[6]), .data5 (in_5[12]), .sel6 (ctl[5]), .data6
       (in_6[12]), .sel7 (ctl[4]), .data7 (in_7[12]), .sel8 (ctl[3]),
       .data8 (in_8[12]), .sel9 (ctl[2]), .data9 (in_9[12]), .sel10
       (ctl[1]), .data10 (in_10[12]), .sel11 (ctl[0]), .data11
       (in_11[12]), .z (z[12]));
  CDN_mux12 g20(.sel0 (ctl[11]), .data0 (in_0[11]), .sel1 (ctl[10]),
       .data1 (in_1[11]), .sel2 (ctl[9]), .data2 (in_2[11]), .sel3
       (ctl[8]), .data3 (in_3[11]), .sel4 (ctl[7]), .data4 (in_4[11]),
       .sel5 (ctl[6]), .data5 (in_5[11]), .sel6 (ctl[5]), .data6
       (in_6[11]), .sel7 (ctl[4]), .data7 (in_7[11]), .sel8 (ctl[3]),
       .data8 (in_8[11]), .sel9 (ctl[2]), .data9 (in_9[11]), .sel10
       (ctl[1]), .data10 (in_10[11]), .sel11 (ctl[0]), .data11
       (in_11[11]), .z (z[11]));
  CDN_mux12 g21(.sel0 (ctl[11]), .data0 (in_0[10]), .sel1 (ctl[10]),
       .data1 (in_1[10]), .sel2 (ctl[9]), .data2 (in_2[10]), .sel3
       (ctl[8]), .data3 (in_3[10]), .sel4 (ctl[7]), .data4 (in_4[10]),
       .sel5 (ctl[6]), .data5 (in_5[10]), .sel6 (ctl[5]), .data6
       (in_6[10]), .sel7 (ctl[4]), .data7 (in_7[10]), .sel8 (ctl[3]),
       .data8 (in_8[10]), .sel9 (ctl[2]), .data9 (in_9[10]), .sel10
       (ctl[1]), .data10 (in_10[10]), .sel11 (ctl[0]), .data11
       (in_11[10]), .z (z[10]));
  CDN_mux12 g22(.sel0 (ctl[11]), .data0 (in_0[9]), .sel1 (ctl[10]),
       .data1 (in_1[9]), .sel2 (ctl[9]), .data2 (in_2[9]), .sel3
       (ctl[8]), .data3 (in_3[9]), .sel4 (ctl[7]), .data4 (in_4[9]),
       .sel5 (ctl[6]), .data5 (in_5[9]), .sel6 (ctl[5]), .data6
       (in_6[9]), .sel7 (ctl[4]), .data7 (in_7[9]), .sel8 (ctl[3]),
       .data8 (in_8[9]), .sel9 (ctl[2]), .data9 (in_9[9]), .sel10
       (ctl[1]), .data10 (in_10[9]), .sel11 (ctl[0]), .data11
       (in_11[9]), .z (z[9]));
  CDN_mux12 g23(.sel0 (ctl[11]), .data0 (in_0[8]), .sel1 (ctl[10]),
       .data1 (in_1[8]), .sel2 (ctl[9]), .data2 (in_2[8]), .sel3
       (ctl[8]), .data3 (in_3[8]), .sel4 (ctl[7]), .data4 (in_4[8]),
       .sel5 (ctl[6]), .data5 (in_5[8]), .sel6 (ctl[5]), .data6
       (in_6[8]), .sel7 (ctl[4]), .data7 (in_7[8]), .sel8 (ctl[3]),
       .data8 (in_8[8]), .sel9 (ctl[2]), .data9 (in_9[8]), .sel10
       (ctl[1]), .data10 (in_10[8]), .sel11 (ctl[0]), .data11
       (in_11[8]), .z (z[8]));
  CDN_mux12 g24(.sel0 (ctl[11]), .data0 (in_0[7]), .sel1 (ctl[10]),
       .data1 (in_1[7]), .sel2 (ctl[9]), .data2 (in_2[7]), .sel3
       (ctl[8]), .data3 (in_3[7]), .sel4 (ctl[7]), .data4 (in_4[7]),
       .sel5 (ctl[6]), .data5 (in_5[7]), .sel6 (ctl[5]), .data6
       (in_6[7]), .sel7 (ctl[4]), .data7 (in_7[7]), .sel8 (ctl[3]),
       .data8 (in_8[7]), .sel9 (ctl[2]), .data9 (in_9[7]), .sel10
       (ctl[1]), .data10 (in_10[7]), .sel11 (ctl[0]), .data11
       (in_11[7]), .z (z[7]));
  CDN_mux12 g25(.sel0 (ctl[11]), .data0 (in_0[6]), .sel1 (ctl[10]),
       .data1 (in_1[6]), .sel2 (ctl[9]), .data2 (in_2[6]), .sel3
       (ctl[8]), .data3 (in_3[6]), .sel4 (ctl[7]), .data4 (in_4[6]),
       .sel5 (ctl[6]), .data5 (in_5[6]), .sel6 (ctl[5]), .data6
       (in_6[6]), .sel7 (ctl[4]), .data7 (in_7[6]), .sel8 (ctl[3]),
       .data8 (in_8[6]), .sel9 (ctl[2]), .data9 (in_9[6]), .sel10
       (ctl[1]), .data10 (in_10[6]), .sel11 (ctl[0]), .data11
       (in_11[6]), .z (z[6]));
  CDN_mux12 g26(.sel0 (ctl[11]), .data0 (in_0[5]), .sel1 (ctl[10]),
       .data1 (in_1[5]), .sel2 (ctl[9]), .data2 (in_2[5]), .sel3
       (ctl[8]), .data3 (in_3[5]), .sel4 (ctl[7]), .data4 (in_4[5]),
       .sel5 (ctl[6]), .data5 (in_5[5]), .sel6 (ctl[5]), .data6
       (in_6[5]), .sel7 (ctl[4]), .data7 (in_7[5]), .sel8 (ctl[3]),
       .data8 (in_8[5]), .sel9 (ctl[2]), .data9 (in_9[5]), .sel10
       (ctl[1]), .data10 (in_10[5]), .sel11 (ctl[0]), .data11
       (in_11[5]), .z (z[5]));
  CDN_mux12 g27(.sel0 (ctl[11]), .data0 (in_0[4]), .sel1 (ctl[10]),
       .data1 (in_1[4]), .sel2 (ctl[9]), .data2 (in_2[4]), .sel3
       (ctl[8]), .data3 (in_3[4]), .sel4 (ctl[7]), .data4 (in_4[4]),
       .sel5 (ctl[6]), .data5 (in_5[4]), .sel6 (ctl[5]), .data6
       (in_6[4]), .sel7 (ctl[4]), .data7 (in_7[4]), .sel8 (ctl[3]),
       .data8 (in_8[4]), .sel9 (ctl[2]), .data9 (in_9[4]), .sel10
       (ctl[1]), .data10 (in_10[4]), .sel11 (ctl[0]), .data11
       (in_11[4]), .z (z[4]));
  CDN_mux12 g28(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g29(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g30(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g31(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_case_box_113(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_116(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_454(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input [12:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  output [12:0] z;
  wire [11:0] ctl;
  wire [12:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  wire [12:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[12]), .sel1 (ctl[10]),
       .data1 (in_1[12]), .sel2 (ctl[9]), .data2 (in_2[12]), .sel3
       (ctl[8]), .data3 (in_3[12]), .sel4 (ctl[7]), .data4 (in_4[12]),
       .sel5 (ctl[6]), .data5 (in_5[12]), .sel6 (ctl[5]), .data6
       (in_6[12]), .sel7 (ctl[4]), .data7 (in_7[12]), .sel8 (ctl[3]),
       .data8 (in_8[12]), .sel9 (ctl[2]), .data9 (in_9[12]), .sel10
       (ctl[1]), .data10 (in_10[12]), .sel11 (ctl[0]), .data11
       (in_11[12]), .z (z[12]));
  CDN_mux12 g14(.sel0 (ctl[11]), .data0 (in_0[11]), .sel1 (ctl[10]),
       .data1 (in_1[11]), .sel2 (ctl[9]), .data2 (in_2[11]), .sel3
       (ctl[8]), .data3 (in_3[11]), .sel4 (ctl[7]), .data4 (in_4[11]),
       .sel5 (ctl[6]), .data5 (in_5[11]), .sel6 (ctl[5]), .data6
       (in_6[11]), .sel7 (ctl[4]), .data7 (in_7[11]), .sel8 (ctl[3]),
       .data8 (in_8[11]), .sel9 (ctl[2]), .data9 (in_9[11]), .sel10
       (ctl[1]), .data10 (in_10[11]), .sel11 (ctl[0]), .data11
       (in_11[11]), .z (z[11]));
  CDN_mux12 g15(.sel0 (ctl[11]), .data0 (in_0[10]), .sel1 (ctl[10]),
       .data1 (in_1[10]), .sel2 (ctl[9]), .data2 (in_2[10]), .sel3
       (ctl[8]), .data3 (in_3[10]), .sel4 (ctl[7]), .data4 (in_4[10]),
       .sel5 (ctl[6]), .data5 (in_5[10]), .sel6 (ctl[5]), .data6
       (in_6[10]), .sel7 (ctl[4]), .data7 (in_7[10]), .sel8 (ctl[3]),
       .data8 (in_8[10]), .sel9 (ctl[2]), .data9 (in_9[10]), .sel10
       (ctl[1]), .data10 (in_10[10]), .sel11 (ctl[0]), .data11
       (in_11[10]), .z (z[10]));
  CDN_mux12 g16(.sel0 (ctl[11]), .data0 (in_0[9]), .sel1 (ctl[10]),
       .data1 (in_1[9]), .sel2 (ctl[9]), .data2 (in_2[9]), .sel3
       (ctl[8]), .data3 (in_3[9]), .sel4 (ctl[7]), .data4 (in_4[9]),
       .sel5 (ctl[6]), .data5 (in_5[9]), .sel6 (ctl[5]), .data6
       (in_6[9]), .sel7 (ctl[4]), .data7 (in_7[9]), .sel8 (ctl[3]),
       .data8 (in_8[9]), .sel9 (ctl[2]), .data9 (in_9[9]), .sel10
       (ctl[1]), .data10 (in_10[9]), .sel11 (ctl[0]), .data11
       (in_11[9]), .z (z[9]));
  CDN_mux12 g17(.sel0 (ctl[11]), .data0 (in_0[8]), .sel1 (ctl[10]),
       .data1 (in_1[8]), .sel2 (ctl[9]), .data2 (in_2[8]), .sel3
       (ctl[8]), .data3 (in_3[8]), .sel4 (ctl[7]), .data4 (in_4[8]),
       .sel5 (ctl[6]), .data5 (in_5[8]), .sel6 (ctl[5]), .data6
       (in_6[8]), .sel7 (ctl[4]), .data7 (in_7[8]), .sel8 (ctl[3]),
       .data8 (in_8[8]), .sel9 (ctl[2]), .data9 (in_9[8]), .sel10
       (ctl[1]), .data10 (in_10[8]), .sel11 (ctl[0]), .data11
       (in_11[8]), .z (z[8]));
  CDN_mux12 g18(.sel0 (ctl[11]), .data0 (in_0[7]), .sel1 (ctl[10]),
       .data1 (in_1[7]), .sel2 (ctl[9]), .data2 (in_2[7]), .sel3
       (ctl[8]), .data3 (in_3[7]), .sel4 (ctl[7]), .data4 (in_4[7]),
       .sel5 (ctl[6]), .data5 (in_5[7]), .sel6 (ctl[5]), .data6
       (in_6[7]), .sel7 (ctl[4]), .data7 (in_7[7]), .sel8 (ctl[3]),
       .data8 (in_8[7]), .sel9 (ctl[2]), .data9 (in_9[7]), .sel10
       (ctl[1]), .data10 (in_10[7]), .sel11 (ctl[0]), .data11
       (in_11[7]), .z (z[7]));
  CDN_mux12 g19(.sel0 (ctl[11]), .data0 (in_0[6]), .sel1 (ctl[10]),
       .data1 (in_1[6]), .sel2 (ctl[9]), .data2 (in_2[6]), .sel3
       (ctl[8]), .data3 (in_3[6]), .sel4 (ctl[7]), .data4 (in_4[6]),
       .sel5 (ctl[6]), .data5 (in_5[6]), .sel6 (ctl[5]), .data6
       (in_6[6]), .sel7 (ctl[4]), .data7 (in_7[6]), .sel8 (ctl[3]),
       .data8 (in_8[6]), .sel9 (ctl[2]), .data9 (in_9[6]), .sel10
       (ctl[1]), .data10 (in_10[6]), .sel11 (ctl[0]), .data11
       (in_11[6]), .z (z[6]));
  CDN_mux12 g20(.sel0 (ctl[11]), .data0 (in_0[5]), .sel1 (ctl[10]),
       .data1 (in_1[5]), .sel2 (ctl[9]), .data2 (in_2[5]), .sel3
       (ctl[8]), .data3 (in_3[5]), .sel4 (ctl[7]), .data4 (in_4[5]),
       .sel5 (ctl[6]), .data5 (in_5[5]), .sel6 (ctl[5]), .data6
       (in_6[5]), .sel7 (ctl[4]), .data7 (in_7[5]), .sel8 (ctl[3]),
       .data8 (in_8[5]), .sel9 (ctl[2]), .data9 (in_9[5]), .sel10
       (ctl[1]), .data10 (in_10[5]), .sel11 (ctl[0]), .data11
       (in_11[5]), .z (z[5]));
  CDN_mux12 g21(.sel0 (ctl[11]), .data0 (in_0[4]), .sel1 (ctl[10]),
       .data1 (in_1[4]), .sel2 (ctl[9]), .data2 (in_2[4]), .sel3
       (ctl[8]), .data3 (in_3[4]), .sel4 (ctl[7]), .data4 (in_4[4]),
       .sel5 (ctl[6]), .data5 (in_5[4]), .sel6 (ctl[5]), .data6
       (in_6[4]), .sel7 (ctl[4]), .data7 (in_7[4]), .sel8 (ctl[3]),
       .data8 (in_8[4]), .sel9 (ctl[2]), .data9 (in_9[4]), .sel10
       (ctl[1]), .data10 (in_10[4]), .sel11 (ctl[0]), .data11
       (in_11[4]), .z (z[4]));
  CDN_mux12 g22(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g23(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g24(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g25(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_case_box_119(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_122(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_125(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_128(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_131(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_520(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input [13:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  output [13:0] z;
  wire [11:0] ctl;
  wire [13:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  wire [13:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[13]), .sel1 (ctl[10]),
       .data1 (in_1[13]), .sel2 (ctl[9]), .data2 (in_2[13]), .sel3
       (ctl[8]), .data3 (in_3[13]), .sel4 (ctl[7]), .data4 (in_4[13]),
       .sel5 (ctl[6]), .data5 (in_5[13]), .sel6 (ctl[5]), .data6
       (in_6[13]), .sel7 (ctl[4]), .data7 (in_7[13]), .sel8 (ctl[3]),
       .data8 (in_8[13]), .sel9 (ctl[2]), .data9 (in_9[13]), .sel10
       (ctl[1]), .data10 (in_10[13]), .sel11 (ctl[0]), .data11
       (in_11[13]), .z (z[13]));
  CDN_mux12 g15(.sel0 (ctl[11]), .data0 (in_0[12]), .sel1 (ctl[10]),
       .data1 (in_1[12]), .sel2 (ctl[9]), .data2 (in_2[12]), .sel3
       (ctl[8]), .data3 (in_3[12]), .sel4 (ctl[7]), .data4 (in_4[12]),
       .sel5 (ctl[6]), .data5 (in_5[12]), .sel6 (ctl[5]), .data6
       (in_6[12]), .sel7 (ctl[4]), .data7 (in_7[12]), .sel8 (ctl[3]),
       .data8 (in_8[12]), .sel9 (ctl[2]), .data9 (in_9[12]), .sel10
       (ctl[1]), .data10 (in_10[12]), .sel11 (ctl[0]), .data11
       (in_11[12]), .z (z[12]));
  CDN_mux12 g16(.sel0 (ctl[11]), .data0 (in_0[11]), .sel1 (ctl[10]),
       .data1 (in_1[11]), .sel2 (ctl[9]), .data2 (in_2[11]), .sel3
       (ctl[8]), .data3 (in_3[11]), .sel4 (ctl[7]), .data4 (in_4[11]),
       .sel5 (ctl[6]), .data5 (in_5[11]), .sel6 (ctl[5]), .data6
       (in_6[11]), .sel7 (ctl[4]), .data7 (in_7[11]), .sel8 (ctl[3]),
       .data8 (in_8[11]), .sel9 (ctl[2]), .data9 (in_9[11]), .sel10
       (ctl[1]), .data10 (in_10[11]), .sel11 (ctl[0]), .data11
       (in_11[11]), .z (z[11]));
  CDN_mux12 g17(.sel0 (ctl[11]), .data0 (in_0[10]), .sel1 (ctl[10]),
       .data1 (in_1[10]), .sel2 (ctl[9]), .data2 (in_2[10]), .sel3
       (ctl[8]), .data3 (in_3[10]), .sel4 (ctl[7]), .data4 (in_4[10]),
       .sel5 (ctl[6]), .data5 (in_5[10]), .sel6 (ctl[5]), .data6
       (in_6[10]), .sel7 (ctl[4]), .data7 (in_7[10]), .sel8 (ctl[3]),
       .data8 (in_8[10]), .sel9 (ctl[2]), .data9 (in_9[10]), .sel10
       (ctl[1]), .data10 (in_10[10]), .sel11 (ctl[0]), .data11
       (in_11[10]), .z (z[10]));
  CDN_mux12 g18(.sel0 (ctl[11]), .data0 (in_0[9]), .sel1 (ctl[10]),
       .data1 (in_1[9]), .sel2 (ctl[9]), .data2 (in_2[9]), .sel3
       (ctl[8]), .data3 (in_3[9]), .sel4 (ctl[7]), .data4 (in_4[9]),
       .sel5 (ctl[6]), .data5 (in_5[9]), .sel6 (ctl[5]), .data6
       (in_6[9]), .sel7 (ctl[4]), .data7 (in_7[9]), .sel8 (ctl[3]),
       .data8 (in_8[9]), .sel9 (ctl[2]), .data9 (in_9[9]), .sel10
       (ctl[1]), .data10 (in_10[9]), .sel11 (ctl[0]), .data11
       (in_11[9]), .z (z[9]));
  CDN_mux12 g19(.sel0 (ctl[11]), .data0 (in_0[8]), .sel1 (ctl[10]),
       .data1 (in_1[8]), .sel2 (ctl[9]), .data2 (in_2[8]), .sel3
       (ctl[8]), .data3 (in_3[8]), .sel4 (ctl[7]), .data4 (in_4[8]),
       .sel5 (ctl[6]), .data5 (in_5[8]), .sel6 (ctl[5]), .data6
       (in_6[8]), .sel7 (ctl[4]), .data7 (in_7[8]), .sel8 (ctl[3]),
       .data8 (in_8[8]), .sel9 (ctl[2]), .data9 (in_9[8]), .sel10
       (ctl[1]), .data10 (in_10[8]), .sel11 (ctl[0]), .data11
       (in_11[8]), .z (z[8]));
  CDN_mux12 g20(.sel0 (ctl[11]), .data0 (in_0[7]), .sel1 (ctl[10]),
       .data1 (in_1[7]), .sel2 (ctl[9]), .data2 (in_2[7]), .sel3
       (ctl[8]), .data3 (in_3[7]), .sel4 (ctl[7]), .data4 (in_4[7]),
       .sel5 (ctl[6]), .data5 (in_5[7]), .sel6 (ctl[5]), .data6
       (in_6[7]), .sel7 (ctl[4]), .data7 (in_7[7]), .sel8 (ctl[3]),
       .data8 (in_8[7]), .sel9 (ctl[2]), .data9 (in_9[7]), .sel10
       (ctl[1]), .data10 (in_10[7]), .sel11 (ctl[0]), .data11
       (in_11[7]), .z (z[7]));
  CDN_mux12 g21(.sel0 (ctl[11]), .data0 (in_0[6]), .sel1 (ctl[10]),
       .data1 (in_1[6]), .sel2 (ctl[9]), .data2 (in_2[6]), .sel3
       (ctl[8]), .data3 (in_3[6]), .sel4 (ctl[7]), .data4 (in_4[6]),
       .sel5 (ctl[6]), .data5 (in_5[6]), .sel6 (ctl[5]), .data6
       (in_6[6]), .sel7 (ctl[4]), .data7 (in_7[6]), .sel8 (ctl[3]),
       .data8 (in_8[6]), .sel9 (ctl[2]), .data9 (in_9[6]), .sel10
       (ctl[1]), .data10 (in_10[6]), .sel11 (ctl[0]), .data11
       (in_11[6]), .z (z[6]));
  CDN_mux12 g22(.sel0 (ctl[11]), .data0 (in_0[5]), .sel1 (ctl[10]),
       .data1 (in_1[5]), .sel2 (ctl[9]), .data2 (in_2[5]), .sel3
       (ctl[8]), .data3 (in_3[5]), .sel4 (ctl[7]), .data4 (in_4[5]),
       .sel5 (ctl[6]), .data5 (in_5[5]), .sel6 (ctl[5]), .data6
       (in_6[5]), .sel7 (ctl[4]), .data7 (in_7[5]), .sel8 (ctl[3]),
       .data8 (in_8[5]), .sel9 (ctl[2]), .data9 (in_9[5]), .sel10
       (ctl[1]), .data10 (in_10[5]), .sel11 (ctl[0]), .data11
       (in_11[5]), .z (z[5]));
  CDN_mux12 g23(.sel0 (ctl[11]), .data0 (in_0[4]), .sel1 (ctl[10]),
       .data1 (in_1[4]), .sel2 (ctl[9]), .data2 (in_2[4]), .sel3
       (ctl[8]), .data3 (in_3[4]), .sel4 (ctl[7]), .data4 (in_4[4]),
       .sel5 (ctl[6]), .data5 (in_5[4]), .sel6 (ctl[5]), .data6
       (in_6[4]), .sel7 (ctl[4]), .data7 (in_7[4]), .sel8 (ctl[3]),
       .data8 (in_8[4]), .sel9 (ctl[2]), .data9 (in_9[4]), .sel10
       (ctl[1]), .data10 (in_10[4]), .sel11 (ctl[0]), .data11
       (in_11[4]), .z (z[4]));
  CDN_mux12 g24(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g25(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g26(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g27(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_case_box_134(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_bmux_546(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, z);
  input [3:0] ctl;
  input [8:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  output [8:0] z;
  wire [3:0] ctl;
  wire [8:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  wire [8:0] z;
  CDN_bmux9 g1(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .sel2
       (ctl[2]), .data4 (in_4[8]), .data5 (in_5[8]), .data6 (in_6[8]),
       .data7 (in_7[8]), .sel3 (ctl[3]), .data8 (in_8[8]), .z (z[8]));
  CDN_bmux9 g2(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .data7 (in_7[7]), .sel3 (ctl[3]), .data8 (in_8[7]), .z (z[7]));
  CDN_bmux9 g3(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .data7 (in_7[6]), .sel3 (ctl[3]), .data8 (in_8[6]), .z (z[6]));
  CDN_bmux9 g4(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .data7 (in_7[5]), .sel3 (ctl[3]), .data8 (in_8[5]), .z (z[5]));
  CDN_bmux9 g5(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .data7 (in_7[4]), .sel3 (ctl[3]), .data8 (in_8[4]), .z (z[4]));
  CDN_bmux9 g6(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .sel3 (ctl[3]), .data8 (in_8[3]), .z (z[3]));
  CDN_bmux9 g7(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .sel3 (ctl[3]), .data8 (in_8[2]), .z (z[2]));
  CDN_bmux9 g8(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .sel3 (ctl[3]), .data8 (in_8[1]), .z (z[1]));
  CDN_bmux9 g9(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .sel3 (ctl[3]), .data8 (in_8[0]), .z (z[0]));
endmodule

module fx68k_case_box_137(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_547(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input [16:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  output [16:0] z;
  wire [11:0] ctl;
  wire [16:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  wire [16:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[16]), .sel1 (ctl[10]),
       .data1 (in_1[16]), .sel2 (ctl[9]), .data2 (in_2[16]), .sel3
       (ctl[8]), .data3 (in_3[16]), .sel4 (ctl[7]), .data4 (in_4[16]),
       .sel5 (ctl[6]), .data5 (in_5[16]), .sel6 (ctl[5]), .data6
       (in_6[16]), .sel7 (ctl[4]), .data7 (in_7[16]), .sel8 (ctl[3]),
       .data8 (in_8[16]), .sel9 (ctl[2]), .data9 (in_9[16]), .sel10
       (ctl[1]), .data10 (in_10[16]), .sel11 (ctl[0]), .data11
       (in_11[16]), .z (z[16]));
  CDN_mux12 g18(.sel0 (ctl[11]), .data0 (in_0[15]), .sel1 (ctl[10]),
       .data1 (in_1[15]), .sel2 (ctl[9]), .data2 (in_2[15]), .sel3
       (ctl[8]), .data3 (in_3[15]), .sel4 (ctl[7]), .data4 (in_4[15]),
       .sel5 (ctl[6]), .data5 (in_5[15]), .sel6 (ctl[5]), .data6
       (in_6[15]), .sel7 (ctl[4]), .data7 (in_7[15]), .sel8 (ctl[3]),
       .data8 (in_8[15]), .sel9 (ctl[2]), .data9 (in_9[15]), .sel10
       (ctl[1]), .data10 (in_10[15]), .sel11 (ctl[0]), .data11
       (in_11[15]), .z (z[15]));
  CDN_mux12 g19(.sel0 (ctl[11]), .data0 (in_0[14]), .sel1 (ctl[10]),
       .data1 (in_1[14]), .sel2 (ctl[9]), .data2 (in_2[14]), .sel3
       (ctl[8]), .data3 (in_3[14]), .sel4 (ctl[7]), .data4 (in_4[14]),
       .sel5 (ctl[6]), .data5 (in_5[14]), .sel6 (ctl[5]), .data6
       (in_6[14]), .sel7 (ctl[4]), .data7 (in_7[14]), .sel8 (ctl[3]),
       .data8 (in_8[14]), .sel9 (ctl[2]), .data9 (in_9[14]), .sel10
       (ctl[1]), .data10 (in_10[14]), .sel11 (ctl[0]), .data11
       (in_11[14]), .z (z[14]));
  CDN_mux12 g20(.sel0 (ctl[11]), .data0 (in_0[13]), .sel1 (ctl[10]),
       .data1 (in_1[13]), .sel2 (ctl[9]), .data2 (in_2[13]), .sel3
       (ctl[8]), .data3 (in_3[13]), .sel4 (ctl[7]), .data4 (in_4[13]),
       .sel5 (ctl[6]), .data5 (in_5[13]), .sel6 (ctl[5]), .data6
       (in_6[13]), .sel7 (ctl[4]), .data7 (in_7[13]), .sel8 (ctl[3]),
       .data8 (in_8[13]), .sel9 (ctl[2]), .data9 (in_9[13]), .sel10
       (ctl[1]), .data10 (in_10[13]), .sel11 (ctl[0]), .data11
       (in_11[13]), .z (z[13]));
  CDN_mux12 g21(.sel0 (ctl[11]), .data0 (in_0[12]), .sel1 (ctl[10]),
       .data1 (in_1[12]), .sel2 (ctl[9]), .data2 (in_2[12]), .sel3
       (ctl[8]), .data3 (in_3[12]), .sel4 (ctl[7]), .data4 (in_4[12]),
       .sel5 (ctl[6]), .data5 (in_5[12]), .sel6 (ctl[5]), .data6
       (in_6[12]), .sel7 (ctl[4]), .data7 (in_7[12]), .sel8 (ctl[3]),
       .data8 (in_8[12]), .sel9 (ctl[2]), .data9 (in_9[12]), .sel10
       (ctl[1]), .data10 (in_10[12]), .sel11 (ctl[0]), .data11
       (in_11[12]), .z (z[12]));
  CDN_mux12 g22(.sel0 (ctl[11]), .data0 (in_0[11]), .sel1 (ctl[10]),
       .data1 (in_1[11]), .sel2 (ctl[9]), .data2 (in_2[11]), .sel3
       (ctl[8]), .data3 (in_3[11]), .sel4 (ctl[7]), .data4 (in_4[11]),
       .sel5 (ctl[6]), .data5 (in_5[11]), .sel6 (ctl[5]), .data6
       (in_6[11]), .sel7 (ctl[4]), .data7 (in_7[11]), .sel8 (ctl[3]),
       .data8 (in_8[11]), .sel9 (ctl[2]), .data9 (in_9[11]), .sel10
       (ctl[1]), .data10 (in_10[11]), .sel11 (ctl[0]), .data11
       (in_11[11]), .z (z[11]));
  CDN_mux12 g23(.sel0 (ctl[11]), .data0 (in_0[10]), .sel1 (ctl[10]),
       .data1 (in_1[10]), .sel2 (ctl[9]), .data2 (in_2[10]), .sel3
       (ctl[8]), .data3 (in_3[10]), .sel4 (ctl[7]), .data4 (in_4[10]),
       .sel5 (ctl[6]), .data5 (in_5[10]), .sel6 (ctl[5]), .data6
       (in_6[10]), .sel7 (ctl[4]), .data7 (in_7[10]), .sel8 (ctl[3]),
       .data8 (in_8[10]), .sel9 (ctl[2]), .data9 (in_9[10]), .sel10
       (ctl[1]), .data10 (in_10[10]), .sel11 (ctl[0]), .data11
       (in_11[10]), .z (z[10]));
  CDN_mux12 g24(.sel0 (ctl[11]), .data0 (in_0[9]), .sel1 (ctl[10]),
       .data1 (in_1[9]), .sel2 (ctl[9]), .data2 (in_2[9]), .sel3
       (ctl[8]), .data3 (in_3[9]), .sel4 (ctl[7]), .data4 (in_4[9]),
       .sel5 (ctl[6]), .data5 (in_5[9]), .sel6 (ctl[5]), .data6
       (in_6[9]), .sel7 (ctl[4]), .data7 (in_7[9]), .sel8 (ctl[3]),
       .data8 (in_8[9]), .sel9 (ctl[2]), .data9 (in_9[9]), .sel10
       (ctl[1]), .data10 (in_10[9]), .sel11 (ctl[0]), .data11
       (in_11[9]), .z (z[9]));
  CDN_mux12 g25(.sel0 (ctl[11]), .data0 (in_0[8]), .sel1 (ctl[10]),
       .data1 (in_1[8]), .sel2 (ctl[9]), .data2 (in_2[8]), .sel3
       (ctl[8]), .data3 (in_3[8]), .sel4 (ctl[7]), .data4 (in_4[8]),
       .sel5 (ctl[6]), .data5 (in_5[8]), .sel6 (ctl[5]), .data6
       (in_6[8]), .sel7 (ctl[4]), .data7 (in_7[8]), .sel8 (ctl[3]),
       .data8 (in_8[8]), .sel9 (ctl[2]), .data9 (in_9[8]), .sel10
       (ctl[1]), .data10 (in_10[8]), .sel11 (ctl[0]), .data11
       (in_11[8]), .z (z[8]));
  CDN_mux12 g26(.sel0 (ctl[11]), .data0 (in_0[7]), .sel1 (ctl[10]),
       .data1 (in_1[7]), .sel2 (ctl[9]), .data2 (in_2[7]), .sel3
       (ctl[8]), .data3 (in_3[7]), .sel4 (ctl[7]), .data4 (in_4[7]),
       .sel5 (ctl[6]), .data5 (in_5[7]), .sel6 (ctl[5]), .data6
       (in_6[7]), .sel7 (ctl[4]), .data7 (in_7[7]), .sel8 (ctl[3]),
       .data8 (in_8[7]), .sel9 (ctl[2]), .data9 (in_9[7]), .sel10
       (ctl[1]), .data10 (in_10[7]), .sel11 (ctl[0]), .data11
       (in_11[7]), .z (z[7]));
  CDN_mux12 g27(.sel0 (ctl[11]), .data0 (in_0[6]), .sel1 (ctl[10]),
       .data1 (in_1[6]), .sel2 (ctl[9]), .data2 (in_2[6]), .sel3
       (ctl[8]), .data3 (in_3[6]), .sel4 (ctl[7]), .data4 (in_4[6]),
       .sel5 (ctl[6]), .data5 (in_5[6]), .sel6 (ctl[5]), .data6
       (in_6[6]), .sel7 (ctl[4]), .data7 (in_7[6]), .sel8 (ctl[3]),
       .data8 (in_8[6]), .sel9 (ctl[2]), .data9 (in_9[6]), .sel10
       (ctl[1]), .data10 (in_10[6]), .sel11 (ctl[0]), .data11
       (in_11[6]), .z (z[6]));
  CDN_mux12 g28(.sel0 (ctl[11]), .data0 (in_0[5]), .sel1 (ctl[10]),
       .data1 (in_1[5]), .sel2 (ctl[9]), .data2 (in_2[5]), .sel3
       (ctl[8]), .data3 (in_3[5]), .sel4 (ctl[7]), .data4 (in_4[5]),
       .sel5 (ctl[6]), .data5 (in_5[5]), .sel6 (ctl[5]), .data6
       (in_6[5]), .sel7 (ctl[4]), .data7 (in_7[5]), .sel8 (ctl[3]),
       .data8 (in_8[5]), .sel9 (ctl[2]), .data9 (in_9[5]), .sel10
       (ctl[1]), .data10 (in_10[5]), .sel11 (ctl[0]), .data11
       (in_11[5]), .z (z[5]));
  CDN_mux12 g29(.sel0 (ctl[11]), .data0 (in_0[4]), .sel1 (ctl[10]),
       .data1 (in_1[4]), .sel2 (ctl[9]), .data2 (in_2[4]), .sel3
       (ctl[8]), .data3 (in_3[4]), .sel4 (ctl[7]), .data4 (in_4[4]),
       .sel5 (ctl[6]), .data5 (in_5[4]), .sel6 (ctl[5]), .data6
       (in_6[4]), .sel7 (ctl[4]), .data7 (in_7[4]), .sel8 (ctl[3]),
       .data8 (in_8[4]), .sel9 (ctl[2]), .data9 (in_9[4]), .sel10
       (ctl[1]), .data10 (in_10[4]), .sel11 (ctl[0]), .data11
       (in_11[4]), .z (z[4]));
  CDN_mux12 g30(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g31(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g32(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g33(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_case_box_140(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_143(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_146(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_149(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_152(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_155(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_158(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_161(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_671(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, z);
  input [8:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  output z;
  wire [8:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  wire z;
  CDN_mux9 g1(.sel0 (ctl[8]), .data0 (in_0), .sel1 (ctl[7]), .data1
       (in_1), .sel2 (ctl[6]), .data2 (in_2), .sel3 (ctl[5]), .data3
       (in_3), .sel4 (ctl[4]), .data4 (in_4), .sel5 (ctl[3]), .data5
       (in_5), .sel6 (ctl[2]), .data6 (in_6), .sel7 (ctl[1]), .data7
       (in_7), .sel8 (ctl[0]), .data8 (in_8), .z (z));
endmodule

module fx68k_case_box_167(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_170(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_173(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_176(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_179(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_182(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_185(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_188(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_191(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_194(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_197(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_200(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_778(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [15:0] z;
  wire [7:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [15:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[15]), .sel1 (ctl[6]), .data1
       (in_1[15]), .sel2 (ctl[5]), .data2 (in_2[15]), .sel3 (ctl[4]),
       .data3 (in_3[15]), .sel4 (ctl[3]), .data4 (in_4[15]), .sel5
       (ctl[2]), .data5 (in_5[15]), .sel6 (ctl[1]), .data6 (in_6[15]),
       .sel7 (ctl[0]), .data7 (in_7[15]), .z (z[15]));
  CDN_mux8 g17(.sel0 (ctl[7]), .data0 (in_0[14]), .sel1 (ctl[6]),
       .data1 (in_1[14]), .sel2 (ctl[5]), .data2 (in_2[14]), .sel3
       (ctl[4]), .data3 (in_3[14]), .sel4 (ctl[3]), .data4 (in_4[14]),
       .sel5 (ctl[2]), .data5 (in_5[14]), .sel6 (ctl[1]), .data6
       (in_6[14]), .sel7 (ctl[0]), .data7 (in_7[14]), .z (z[14]));
  CDN_mux8 g18(.sel0 (ctl[7]), .data0 (in_0[13]), .sel1 (ctl[6]),
       .data1 (in_1[13]), .sel2 (ctl[5]), .data2 (in_2[13]), .sel3
       (ctl[4]), .data3 (in_3[13]), .sel4 (ctl[3]), .data4 (in_4[13]),
       .sel5 (ctl[2]), .data5 (in_5[13]), .sel6 (ctl[1]), .data6
       (in_6[13]), .sel7 (ctl[0]), .data7 (in_7[13]), .z (z[13]));
  CDN_mux8 g19(.sel0 (ctl[7]), .data0 (in_0[12]), .sel1 (ctl[6]),
       .data1 (in_1[12]), .sel2 (ctl[5]), .data2 (in_2[12]), .sel3
       (ctl[4]), .data3 (in_3[12]), .sel4 (ctl[3]), .data4 (in_4[12]),
       .sel5 (ctl[2]), .data5 (in_5[12]), .sel6 (ctl[1]), .data6
       (in_6[12]), .sel7 (ctl[0]), .data7 (in_7[12]), .z (z[12]));
  CDN_mux8 g20(.sel0 (ctl[7]), .data0 (in_0[11]), .sel1 (ctl[6]),
       .data1 (in_1[11]), .sel2 (ctl[5]), .data2 (in_2[11]), .sel3
       (ctl[4]), .data3 (in_3[11]), .sel4 (ctl[3]), .data4 (in_4[11]),
       .sel5 (ctl[2]), .data5 (in_5[11]), .sel6 (ctl[1]), .data6
       (in_6[11]), .sel7 (ctl[0]), .data7 (in_7[11]), .z (z[11]));
  CDN_mux8 g21(.sel0 (ctl[7]), .data0 (in_0[10]), .sel1 (ctl[6]),
       .data1 (in_1[10]), .sel2 (ctl[5]), .data2 (in_2[10]), .sel3
       (ctl[4]), .data3 (in_3[10]), .sel4 (ctl[3]), .data4 (in_4[10]),
       .sel5 (ctl[2]), .data5 (in_5[10]), .sel6 (ctl[1]), .data6
       (in_6[10]), .sel7 (ctl[0]), .data7 (in_7[10]), .z (z[10]));
  CDN_mux8 g22(.sel0 (ctl[7]), .data0 (in_0[9]), .sel1 (ctl[6]), .data1
       (in_1[9]), .sel2 (ctl[5]), .data2 (in_2[9]), .sel3 (ctl[4]),
       .data3 (in_3[9]), .sel4 (ctl[3]), .data4 (in_4[9]), .sel5
       (ctl[2]), .data5 (in_5[9]), .sel6 (ctl[1]), .data6 (in_6[9]),
       .sel7 (ctl[0]), .data7 (in_7[9]), .z (z[9]));
  CDN_mux8 g23(.sel0 (ctl[7]), .data0 (in_0[8]), .sel1 (ctl[6]), .data1
       (in_1[8]), .sel2 (ctl[5]), .data2 (in_2[8]), .sel3 (ctl[4]),
       .data3 (in_3[8]), .sel4 (ctl[3]), .data4 (in_4[8]), .sel5
       (ctl[2]), .data5 (in_5[8]), .sel6 (ctl[1]), .data6 (in_6[8]),
       .sel7 (ctl[0]), .data7 (in_7[8]), .z (z[8]));
  CDN_mux8 g24(.sel0 (ctl[7]), .data0 (in_0[7]), .sel1 (ctl[6]), .data1
       (in_1[7]), .sel2 (ctl[5]), .data2 (in_2[7]), .sel3 (ctl[4]),
       .data3 (in_3[7]), .sel4 (ctl[3]), .data4 (in_4[7]), .sel5
       (ctl[2]), .data5 (in_5[7]), .sel6 (ctl[1]), .data6 (in_6[7]),
       .sel7 (ctl[0]), .data7 (in_7[7]), .z (z[7]));
  CDN_mux8 g25(.sel0 (ctl[7]), .data0 (in_0[6]), .sel1 (ctl[6]), .data1
       (in_1[6]), .sel2 (ctl[5]), .data2 (in_2[6]), .sel3 (ctl[4]),
       .data3 (in_3[6]), .sel4 (ctl[3]), .data4 (in_4[6]), .sel5
       (ctl[2]), .data5 (in_5[6]), .sel6 (ctl[1]), .data6 (in_6[6]),
       .sel7 (ctl[0]), .data7 (in_7[6]), .z (z[6]));
  CDN_mux8 g26(.sel0 (ctl[7]), .data0 (in_0[5]), .sel1 (ctl[6]), .data1
       (in_1[5]), .sel2 (ctl[5]), .data2 (in_2[5]), .sel3 (ctl[4]),
       .data3 (in_3[5]), .sel4 (ctl[3]), .data4 (in_4[5]), .sel5
       (ctl[2]), .data5 (in_5[5]), .sel6 (ctl[1]), .data6 (in_6[5]),
       .sel7 (ctl[0]), .data7 (in_7[5]), .z (z[5]));
  CDN_mux8 g27(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g28(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g29(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g30(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g31(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_203(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_793(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, z);
  input [10:0] ctl;
  input [11:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  output [11:0] z;
  wire [10:0] ctl;
  wire [11:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10;
  wire [11:0] z;
  CDN_mux11 g1(.sel0 (ctl[10]), .data0 (in_0[11]), .sel1 (ctl[9]),
       .data1 (in_1[11]), .sel2 (ctl[8]), .data2 (in_2[11]), .sel3
       (ctl[7]), .data3 (in_3[11]), .sel4 (ctl[6]), .data4 (in_4[11]),
       .sel5 (ctl[5]), .data5 (in_5[11]), .sel6 (ctl[4]), .data6
       (in_6[11]), .sel7 (ctl[3]), .data7 (in_7[11]), .sel8 (ctl[2]),
       .data8 (in_8[11]), .sel9 (ctl[1]), .data9 (in_9[11]), .sel10
       (ctl[0]), .data10 (in_10[11]), .z (z[11]));
  CDN_mux11 g13(.sel0 (ctl[10]), .data0 (in_0[10]), .sel1 (ctl[9]),
       .data1 (in_1[10]), .sel2 (ctl[8]), .data2 (in_2[10]), .sel3
       (ctl[7]), .data3 (in_3[10]), .sel4 (ctl[6]), .data4 (in_4[10]),
       .sel5 (ctl[5]), .data5 (in_5[10]), .sel6 (ctl[4]), .data6
       (in_6[10]), .sel7 (ctl[3]), .data7 (in_7[10]), .sel8 (ctl[2]),
       .data8 (in_8[10]), .sel9 (ctl[1]), .data9 (in_9[10]), .sel10
       (ctl[0]), .data10 (in_10[10]), .z (z[10]));
  CDN_mux11 g14(.sel0 (ctl[10]), .data0 (in_0[9]), .sel1 (ctl[9]),
       .data1 (in_1[9]), .sel2 (ctl[8]), .data2 (in_2[9]), .sel3
       (ctl[7]), .data3 (in_3[9]), .sel4 (ctl[6]), .data4 (in_4[9]),
       .sel5 (ctl[5]), .data5 (in_5[9]), .sel6 (ctl[4]), .data6
       (in_6[9]), .sel7 (ctl[3]), .data7 (in_7[9]), .sel8 (ctl[2]),
       .data8 (in_8[9]), .sel9 (ctl[1]), .data9 (in_9[9]), .sel10
       (ctl[0]), .data10 (in_10[9]), .z (z[9]));
  CDN_mux11 g15(.sel0 (ctl[10]), .data0 (in_0[8]), .sel1 (ctl[9]),
       .data1 (in_1[8]), .sel2 (ctl[8]), .data2 (in_2[8]), .sel3
       (ctl[7]), .data3 (in_3[8]), .sel4 (ctl[6]), .data4 (in_4[8]),
       .sel5 (ctl[5]), .data5 (in_5[8]), .sel6 (ctl[4]), .data6
       (in_6[8]), .sel7 (ctl[3]), .data7 (in_7[8]), .sel8 (ctl[2]),
       .data8 (in_8[8]), .sel9 (ctl[1]), .data9 (in_9[8]), .sel10
       (ctl[0]), .data10 (in_10[8]), .z (z[8]));
  CDN_mux11 g16(.sel0 (ctl[10]), .data0 (in_0[7]), .sel1 (ctl[9]),
       .data1 (in_1[7]), .sel2 (ctl[8]), .data2 (in_2[7]), .sel3
       (ctl[7]), .data3 (in_3[7]), .sel4 (ctl[6]), .data4 (in_4[7]),
       .sel5 (ctl[5]), .data5 (in_5[7]), .sel6 (ctl[4]), .data6
       (in_6[7]), .sel7 (ctl[3]), .data7 (in_7[7]), .sel8 (ctl[2]),
       .data8 (in_8[7]), .sel9 (ctl[1]), .data9 (in_9[7]), .sel10
       (ctl[0]), .data10 (in_10[7]), .z (z[7]));
  CDN_mux11 g17(.sel0 (ctl[10]), .data0 (in_0[6]), .sel1 (ctl[9]),
       .data1 (in_1[6]), .sel2 (ctl[8]), .data2 (in_2[6]), .sel3
       (ctl[7]), .data3 (in_3[6]), .sel4 (ctl[6]), .data4 (in_4[6]),
       .sel5 (ctl[5]), .data5 (in_5[6]), .sel6 (ctl[4]), .data6
       (in_6[6]), .sel7 (ctl[3]), .data7 (in_7[6]), .sel8 (ctl[2]),
       .data8 (in_8[6]), .sel9 (ctl[1]), .data9 (in_9[6]), .sel10
       (ctl[0]), .data10 (in_10[6]), .z (z[6]));
  CDN_mux11 g18(.sel0 (ctl[10]), .data0 (in_0[5]), .sel1 (ctl[9]),
       .data1 (in_1[5]), .sel2 (ctl[8]), .data2 (in_2[5]), .sel3
       (ctl[7]), .data3 (in_3[5]), .sel4 (ctl[6]), .data4 (in_4[5]),
       .sel5 (ctl[5]), .data5 (in_5[5]), .sel6 (ctl[4]), .data6
       (in_6[5]), .sel7 (ctl[3]), .data7 (in_7[5]), .sel8 (ctl[2]),
       .data8 (in_8[5]), .sel9 (ctl[1]), .data9 (in_9[5]), .sel10
       (ctl[0]), .data10 (in_10[5]), .z (z[5]));
  CDN_mux11 g19(.sel0 (ctl[10]), .data0 (in_0[4]), .sel1 (ctl[9]),
       .data1 (in_1[4]), .sel2 (ctl[8]), .data2 (in_2[4]), .sel3
       (ctl[7]), .data3 (in_3[4]), .sel4 (ctl[6]), .data4 (in_4[4]),
       .sel5 (ctl[5]), .data5 (in_5[4]), .sel6 (ctl[4]), .data6
       (in_6[4]), .sel7 (ctl[3]), .data7 (in_7[4]), .sel8 (ctl[2]),
       .data8 (in_8[4]), .sel9 (ctl[1]), .data9 (in_9[4]), .sel10
       (ctl[0]), .data10 (in_10[4]), .z (z[4]));
  CDN_mux11 g20(.sel0 (ctl[10]), .data0 (in_0[3]), .sel1 (ctl[9]),
       .data1 (in_1[3]), .sel2 (ctl[8]), .data2 (in_2[3]), .sel3
       (ctl[7]), .data3 (in_3[3]), .sel4 (ctl[6]), .data4 (in_4[3]),
       .sel5 (ctl[5]), .data5 (in_5[3]), .sel6 (ctl[4]), .data6
       (in_6[3]), .sel7 (ctl[3]), .data7 (in_7[3]), .sel8 (ctl[2]),
       .data8 (in_8[3]), .sel9 (ctl[1]), .data9 (in_9[3]), .sel10
       (ctl[0]), .data10 (in_10[3]), .z (z[3]));
  CDN_mux11 g21(.sel0 (ctl[10]), .data0 (in_0[2]), .sel1 (ctl[9]),
       .data1 (in_1[2]), .sel2 (ctl[8]), .data2 (in_2[2]), .sel3
       (ctl[7]), .data3 (in_3[2]), .sel4 (ctl[6]), .data4 (in_4[2]),
       .sel5 (ctl[5]), .data5 (in_5[2]), .sel6 (ctl[4]), .data6
       (in_6[2]), .sel7 (ctl[3]), .data7 (in_7[2]), .sel8 (ctl[2]),
       .data8 (in_8[2]), .sel9 (ctl[1]), .data9 (in_9[2]), .sel10
       (ctl[0]), .data10 (in_10[2]), .z (z[2]));
  CDN_mux11 g22(.sel0 (ctl[10]), .data0 (in_0[1]), .sel1 (ctl[9]),
       .data1 (in_1[1]), .sel2 (ctl[8]), .data2 (in_2[1]), .sel3
       (ctl[7]), .data3 (in_3[1]), .sel4 (ctl[6]), .data4 (in_4[1]),
       .sel5 (ctl[5]), .data5 (in_5[1]), .sel6 (ctl[4]), .data6
       (in_6[1]), .sel7 (ctl[3]), .data7 (in_7[1]), .sel8 (ctl[2]),
       .data8 (in_8[1]), .sel9 (ctl[1]), .data9 (in_9[1]), .sel10
       (ctl[0]), .data10 (in_10[1]), .z (z[1]));
  CDN_mux11 g23(.sel0 (ctl[10]), .data0 (in_0[0]), .sel1 (ctl[9]),
       .data1 (in_1[0]), .sel2 (ctl[8]), .data2 (in_2[0]), .sel3
       (ctl[7]), .data3 (in_3[0]), .sel4 (ctl[6]), .data4 (in_4[0]),
       .sel5 (ctl[5]), .data5 (in_5[0]), .sel6 (ctl[4]), .data6
       (in_6[0]), .sel7 (ctl[3]), .data7 (in_7[0]), .sel8 (ctl[2]),
       .data8 (in_8[0]), .sel9 (ctl[1]), .data9 (in_9[0]), .sel10
       (ctl[0]), .data10 (in_10[0]), .z (z[0]));
endmodule

module fx68k_mux_804(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, z);
  input [8:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  output [8:0] z;
  wire [8:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  wire [8:0] z;
  CDN_mux9 g1(.sel0 (ctl[8]), .data0 (in_0[8]), .sel1 (ctl[7]), .data1
       (in_1[8]), .sel2 (ctl[6]), .data2 (in_2[8]), .sel3 (ctl[5]),
       .data3 (in_3[8]), .sel4 (ctl[4]), .data4 (in_4[8]), .sel5
       (ctl[3]), .data5 (in_5[8]), .sel6 (ctl[2]), .data6 (in_6[8]),
       .sel7 (ctl[1]), .data7 (in_7[8]), .sel8 (ctl[0]), .data8
       (in_8[8]), .z (z[8]));
  CDN_mux9 g10(.sel0 (ctl[8]), .data0 (in_0[7]), .sel1 (ctl[7]), .data1
       (in_1[7]), .sel2 (ctl[6]), .data2 (in_2[7]), .sel3 (ctl[5]),
       .data3 (in_3[7]), .sel4 (ctl[4]), .data4 (in_4[7]), .sel5
       (ctl[3]), .data5 (in_5[7]), .sel6 (ctl[2]), .data6 (in_6[7]),
       .sel7 (ctl[1]), .data7 (in_7[7]), .sel8 (ctl[0]), .data8
       (in_8[7]), .z (z[7]));
  CDN_mux9 g11(.sel0 (ctl[8]), .data0 (in_0[6]), .sel1 (ctl[7]), .data1
       (in_1[6]), .sel2 (ctl[6]), .data2 (in_2[6]), .sel3 (ctl[5]),
       .data3 (in_3[6]), .sel4 (ctl[4]), .data4 (in_4[6]), .sel5
       (ctl[3]), .data5 (in_5[6]), .sel6 (ctl[2]), .data6 (in_6[6]),
       .sel7 (ctl[1]), .data7 (in_7[6]), .sel8 (ctl[0]), .data8
       (in_8[6]), .z (z[6]));
  CDN_mux9 g12(.sel0 (ctl[8]), .data0 (in_0[5]), .sel1 (ctl[7]), .data1
       (in_1[5]), .sel2 (ctl[6]), .data2 (in_2[5]), .sel3 (ctl[5]),
       .data3 (in_3[5]), .sel4 (ctl[4]), .data4 (in_4[5]), .sel5
       (ctl[3]), .data5 (in_5[5]), .sel6 (ctl[2]), .data6 (in_6[5]),
       .sel7 (ctl[1]), .data7 (in_7[5]), .sel8 (ctl[0]), .data8
       (in_8[5]), .z (z[5]));
  CDN_mux9 g13(.sel0 (ctl[8]), .data0 (in_0[4]), .sel1 (ctl[7]), .data1
       (in_1[4]), .sel2 (ctl[6]), .data2 (in_2[4]), .sel3 (ctl[5]),
       .data3 (in_3[4]), .sel4 (ctl[4]), .data4 (in_4[4]), .sel5
       (ctl[3]), .data5 (in_5[4]), .sel6 (ctl[2]), .data6 (in_6[4]),
       .sel7 (ctl[1]), .data7 (in_7[4]), .sel8 (ctl[0]), .data8
       (in_8[4]), .z (z[4]));
  CDN_mux9 g14(.sel0 (ctl[8]), .data0 (in_0[3]), .sel1 (ctl[7]), .data1
       (in_1[3]), .sel2 (ctl[6]), .data2 (in_2[3]), .sel3 (ctl[5]),
       .data3 (in_3[3]), .sel4 (ctl[4]), .data4 (in_4[3]), .sel5
       (ctl[3]), .data5 (in_5[3]), .sel6 (ctl[2]), .data6 (in_6[3]),
       .sel7 (ctl[1]), .data7 (in_7[3]), .sel8 (ctl[0]), .data8
       (in_8[3]), .z (z[3]));
  CDN_mux9 g15(.sel0 (ctl[8]), .data0 (in_0[2]), .sel1 (ctl[7]), .data1
       (in_1[2]), .sel2 (ctl[6]), .data2 (in_2[2]), .sel3 (ctl[5]),
       .data3 (in_3[2]), .sel4 (ctl[4]), .data4 (in_4[2]), .sel5
       (ctl[3]), .data5 (in_5[2]), .sel6 (ctl[2]), .data6 (in_6[2]),
       .sel7 (ctl[1]), .data7 (in_7[2]), .sel8 (ctl[0]), .data8
       (in_8[2]), .z (z[2]));
  CDN_mux9 g16(.sel0 (ctl[8]), .data0 (in_0[1]), .sel1 (ctl[7]), .data1
       (in_1[1]), .sel2 (ctl[6]), .data2 (in_2[1]), .sel3 (ctl[5]),
       .data3 (in_3[1]), .sel4 (ctl[4]), .data4 (in_4[1]), .sel5
       (ctl[3]), .data5 (in_5[1]), .sel6 (ctl[2]), .data6 (in_6[1]),
       .sel7 (ctl[1]), .data7 (in_7[1]), .sel8 (ctl[0]), .data8
       (in_8[1]), .z (z[1]));
  CDN_mux9 g17(.sel0 (ctl[8]), .data0 (in_0[0]), .sel1 (ctl[7]), .data1
       (in_1[0]), .sel2 (ctl[6]), .data2 (in_2[0]), .sel3 (ctl[5]),
       .data3 (in_3[0]), .sel4 (ctl[4]), .data4 (in_4[0]), .sel5
       (ctl[3]), .data5 (in_5[0]), .sel6 (ctl[2]), .data6 (in_6[0]),
       .sel7 (ctl[1]), .data7 (in_7[0]), .sel8 (ctl[0]), .data8
       (in_8[0]), .z (z[0]));
endmodule

module fx68k_mux_812(ctl, in_0, in_1, in_2, in_3, z);
  input [3:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3;
  output [9:0] z;
  wire [3:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3;
  wire [9:0] z;
  CDN_mux4 g1(.sel0 (ctl[3]), .data0 (in_0[9]), .sel1 (ctl[2]), .data1
       (in_1[9]), .sel2 (ctl[1]), .data2 (in_2[9]), .sel3 (ctl[0]),
       .data3 (in_3[9]), .z (z[9]));
  CDN_mux4 g11(.sel0 (ctl[3]), .data0 (in_0[8]), .sel1 (ctl[2]), .data1
       (in_1[8]), .sel2 (ctl[1]), .data2 (in_2[8]), .sel3 (ctl[0]),
       .data3 (in_3[8]), .z (z[8]));
  CDN_mux4 g12(.sel0 (ctl[3]), .data0 (in_0[7]), .sel1 (ctl[2]), .data1
       (in_1[7]), .sel2 (ctl[1]), .data2 (in_2[7]), .sel3 (ctl[0]),
       .data3 (in_3[7]), .z (z[7]));
  CDN_mux4 g13(.sel0 (ctl[3]), .data0 (in_0[6]), .sel1 (ctl[2]), .data1
       (in_1[6]), .sel2 (ctl[1]), .data2 (in_2[6]), .sel3 (ctl[0]),
       .data3 (in_3[6]), .z (z[6]));
  CDN_mux4 g14(.sel0 (ctl[3]), .data0 (in_0[5]), .sel1 (ctl[2]), .data1
       (in_1[5]), .sel2 (ctl[1]), .data2 (in_2[5]), .sel3 (ctl[0]),
       .data3 (in_3[5]), .z (z[5]));
  CDN_mux4 g15(.sel0 (ctl[3]), .data0 (in_0[4]), .sel1 (ctl[2]), .data1
       (in_1[4]), .sel2 (ctl[1]), .data2 (in_2[4]), .sel3 (ctl[0]),
       .data3 (in_3[4]), .z (z[4]));
  CDN_mux4 g16(.sel0 (ctl[3]), .data0 (in_0[3]), .sel1 (ctl[2]), .data1
       (in_1[3]), .sel2 (ctl[1]), .data2 (in_2[3]), .sel3 (ctl[0]),
       .data3 (in_3[3]), .z (z[3]));
  CDN_mux4 g17(.sel0 (ctl[3]), .data0 (in_0[2]), .sel1 (ctl[2]), .data1
       (in_1[2]), .sel2 (ctl[1]), .data2 (in_2[2]), .sel3 (ctl[0]),
       .data3 (in_3[2]), .z (z[2]));
  CDN_mux4 g18(.sel0 (ctl[3]), .data0 (in_0[1]), .sel1 (ctl[2]), .data1
       (in_1[1]), .sel2 (ctl[1]), .data2 (in_2[1]), .sel3 (ctl[0]),
       .data3 (in_3[1]), .z (z[1]));
  CDN_mux4 g19(.sel0 (ctl[3]), .data0 (in_0[0]), .sel1 (ctl[2]), .data1
       (in_1[0]), .sel2 (ctl[1]), .data2 (in_2[0]), .sel3 (ctl[0]),
       .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_case_box_212(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_case_box_215(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_case_box_218(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_case_box_221(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_case_box_224(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_case_box_227(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_case_box_230(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_case_box_233(in_0, out_0);
  input [3:0] in_0;
  output [9:0] out_0;
  wire [3:0] in_0;
  wire [9:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_16, n_18;
  wire n_87, n_88;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[3];
  nor g1 (out_0[9], n_5, n_10);
  nand g2 (n_5, n_87, n_88);
  not g3 (n_87, in_0[3]);
  not g4 (n_88, in_0[0]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[2]);
  not g7 (n_9, in_0[1]);
  nor g8 (out_0[8], in_0[2], n_12);
  nand g9 (n_12, n_9, in_0[0]);
  nor g10 (out_0[7], in_0[2], n_14);
  nand g11 (n_14, in_0[1], n_88);
  nor g12 (out_0[6], in_0[2], n_16);
  nand g13 (n_16, in_0[1], in_0[0]);
  nor g14 (out_0[5], n_7, n_18);
  nand g15 (n_18, n_9, n_88);
  nor g16 (out_0[4], n_12, n_7);
  nor g17 (out_0[3], n_14, n_7);
  nor g18 (out_0[2], n_16, n_7);
endmodule

module fx68k_mux_893(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [6:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [6:0] z;
  wire [7:0] ctl;
  wire [6:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [6:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[6]), .sel1 (ctl[6]), .data1
       (in_1[6]), .sel2 (ctl[5]), .data2 (in_2[6]), .sel3 (ctl[4]),
       .data3 (in_3[6]), .sel4 (ctl[3]), .data4 (in_4[6]), .sel5
       (ctl[2]), .data5 (in_5[6]), .sel6 (ctl[1]), .data6 (in_6[6]),
       .sel7 (ctl[0]), .data7 (in_7[6]), .z (z[6]));
  CDN_mux8 g8(.sel0 (ctl[7]), .data0 (in_0[5]), .sel1 (ctl[6]), .data1
       (in_1[5]), .sel2 (ctl[5]), .data2 (in_2[5]), .sel3 (ctl[4]),
       .data3 (in_3[5]), .sel4 (ctl[3]), .data4 (in_4[5]), .sel5
       (ctl[2]), .data5 (in_5[5]), .sel6 (ctl[1]), .data6 (in_6[5]),
       .sel7 (ctl[0]), .data7 (in_7[5]), .z (z[5]));
  CDN_mux8 g9(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g10(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g11(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g12(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g13(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_239(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_899(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, z);
  input [10:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7,
       in_8, in_9, in_10;
  output [10:0] z;
  wire [10:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7,
       in_8, in_9, in_10;
  wire [10:0] z;
  CDN_mux11 g1(.sel0 (ctl[10]), .data0 (in_0[10]), .sel1 (ctl[9]),
       .data1 (in_1[10]), .sel2 (ctl[8]), .data2 (in_2[10]), .sel3
       (ctl[7]), .data3 (in_3[10]), .sel4 (ctl[6]), .data4 (in_4[10]),
       .sel5 (ctl[5]), .data5 (in_5[10]), .sel6 (ctl[4]), .data6
       (in_6[10]), .sel7 (ctl[3]), .data7 (in_7[10]), .sel8 (ctl[2]),
       .data8 (in_8[10]), .sel9 (ctl[1]), .data9 (in_9[10]), .sel10
       (ctl[0]), .data10 (in_10[10]), .z (z[10]));
  CDN_mux11 g12(.sel0 (ctl[10]), .data0 (in_0[9]), .sel1 (ctl[9]),
       .data1 (in_1[9]), .sel2 (ctl[8]), .data2 (in_2[9]), .sel3
       (ctl[7]), .data3 (in_3[9]), .sel4 (ctl[6]), .data4 (in_4[9]),
       .sel5 (ctl[5]), .data5 (in_5[9]), .sel6 (ctl[4]), .data6
       (in_6[9]), .sel7 (ctl[3]), .data7 (in_7[9]), .sel8 (ctl[2]),
       .data8 (in_8[9]), .sel9 (ctl[1]), .data9 (in_9[9]), .sel10
       (ctl[0]), .data10 (in_10[9]), .z (z[9]));
  CDN_mux11 g13(.sel0 (ctl[10]), .data0 (in_0[8]), .sel1 (ctl[9]),
       .data1 (in_1[8]), .sel2 (ctl[8]), .data2 (in_2[8]), .sel3
       (ctl[7]), .data3 (in_3[8]), .sel4 (ctl[6]), .data4 (in_4[8]),
       .sel5 (ctl[5]), .data5 (in_5[8]), .sel6 (ctl[4]), .data6
       (in_6[8]), .sel7 (ctl[3]), .data7 (in_7[8]), .sel8 (ctl[2]),
       .data8 (in_8[8]), .sel9 (ctl[1]), .data9 (in_9[8]), .sel10
       (ctl[0]), .data10 (in_10[8]), .z (z[8]));
  CDN_mux11 g14(.sel0 (ctl[10]), .data0 (in_0[7]), .sel1 (ctl[9]),
       .data1 (in_1[7]), .sel2 (ctl[8]), .data2 (in_2[7]), .sel3
       (ctl[7]), .data3 (in_3[7]), .sel4 (ctl[6]), .data4 (in_4[7]),
       .sel5 (ctl[5]), .data5 (in_5[7]), .sel6 (ctl[4]), .data6
       (in_6[7]), .sel7 (ctl[3]), .data7 (in_7[7]), .sel8 (ctl[2]),
       .data8 (in_8[7]), .sel9 (ctl[1]), .data9 (in_9[7]), .sel10
       (ctl[0]), .data10 (in_10[7]), .z (z[7]));
  CDN_mux11 g15(.sel0 (ctl[10]), .data0 (in_0[6]), .sel1 (ctl[9]),
       .data1 (in_1[6]), .sel2 (ctl[8]), .data2 (in_2[6]), .sel3
       (ctl[7]), .data3 (in_3[6]), .sel4 (ctl[6]), .data4 (in_4[6]),
       .sel5 (ctl[5]), .data5 (in_5[6]), .sel6 (ctl[4]), .data6
       (in_6[6]), .sel7 (ctl[3]), .data7 (in_7[6]), .sel8 (ctl[2]),
       .data8 (in_8[6]), .sel9 (ctl[1]), .data9 (in_9[6]), .sel10
       (ctl[0]), .data10 (in_10[6]), .z (z[6]));
  CDN_mux11 g16(.sel0 (ctl[10]), .data0 (in_0[5]), .sel1 (ctl[9]),
       .data1 (in_1[5]), .sel2 (ctl[8]), .data2 (in_2[5]), .sel3
       (ctl[7]), .data3 (in_3[5]), .sel4 (ctl[6]), .data4 (in_4[5]),
       .sel5 (ctl[5]), .data5 (in_5[5]), .sel6 (ctl[4]), .data6
       (in_6[5]), .sel7 (ctl[3]), .data7 (in_7[5]), .sel8 (ctl[2]),
       .data8 (in_8[5]), .sel9 (ctl[1]), .data9 (in_9[5]), .sel10
       (ctl[0]), .data10 (in_10[5]), .z (z[5]));
  CDN_mux11 g17(.sel0 (ctl[10]), .data0 (in_0[4]), .sel1 (ctl[9]),
       .data1 (in_1[4]), .sel2 (ctl[8]), .data2 (in_2[4]), .sel3
       (ctl[7]), .data3 (in_3[4]), .sel4 (ctl[6]), .data4 (in_4[4]),
       .sel5 (ctl[5]), .data5 (in_5[4]), .sel6 (ctl[4]), .data6
       (in_6[4]), .sel7 (ctl[3]), .data7 (in_7[4]), .sel8 (ctl[2]),
       .data8 (in_8[4]), .sel9 (ctl[1]), .data9 (in_9[4]), .sel10
       (ctl[0]), .data10 (in_10[4]), .z (z[4]));
  CDN_mux11 g18(.sel0 (ctl[10]), .data0 (in_0[3]), .sel1 (ctl[9]),
       .data1 (in_1[3]), .sel2 (ctl[8]), .data2 (in_2[3]), .sel3
       (ctl[7]), .data3 (in_3[3]), .sel4 (ctl[6]), .data4 (in_4[3]),
       .sel5 (ctl[5]), .data5 (in_5[3]), .sel6 (ctl[4]), .data6
       (in_6[3]), .sel7 (ctl[3]), .data7 (in_7[3]), .sel8 (ctl[2]),
       .data8 (in_8[3]), .sel9 (ctl[1]), .data9 (in_9[3]), .sel10
       (ctl[0]), .data10 (in_10[3]), .z (z[3]));
  CDN_mux11 g19(.sel0 (ctl[10]), .data0 (in_0[2]), .sel1 (ctl[9]),
       .data1 (in_1[2]), .sel2 (ctl[8]), .data2 (in_2[2]), .sel3
       (ctl[7]), .data3 (in_3[2]), .sel4 (ctl[6]), .data4 (in_4[2]),
       .sel5 (ctl[5]), .data5 (in_5[2]), .sel6 (ctl[4]), .data6
       (in_6[2]), .sel7 (ctl[3]), .data7 (in_7[2]), .sel8 (ctl[2]),
       .data8 (in_8[2]), .sel9 (ctl[1]), .data9 (in_9[2]), .sel10
       (ctl[0]), .data10 (in_10[2]), .z (z[2]));
  CDN_mux11 g20(.sel0 (ctl[10]), .data0 (in_0[1]), .sel1 (ctl[9]),
       .data1 (in_1[1]), .sel2 (ctl[8]), .data2 (in_2[1]), .sel3
       (ctl[7]), .data3 (in_3[1]), .sel4 (ctl[6]), .data4 (in_4[1]),
       .sel5 (ctl[5]), .data5 (in_5[1]), .sel6 (ctl[4]), .data6
       (in_6[1]), .sel7 (ctl[3]), .data7 (in_7[1]), .sel8 (ctl[2]),
       .data8 (in_8[1]), .sel9 (ctl[1]), .data9 (in_9[1]), .sel10
       (ctl[0]), .data10 (in_10[1]), .z (z[1]));
  CDN_mux11 g21(.sel0 (ctl[10]), .data0 (in_0[0]), .sel1 (ctl[9]),
       .data1 (in_1[0]), .sel2 (ctl[8]), .data2 (in_2[0]), .sel3
       (ctl[7]), .data3 (in_3[0]), .sel4 (ctl[6]), .data4 (in_4[0]),
       .sel5 (ctl[5]), .data5 (in_5[0]), .sel6 (ctl[4]), .data6
       (in_6[0]), .sel7 (ctl[3]), .data7 (in_7[0]), .sel8 (ctl[2]),
       .data8 (in_8[0]), .sel9 (ctl[1]), .data9 (in_9[0]), .sel10
       (ctl[0]), .data10 (in_10[0]), .z (z[0]));
endmodule

module fx68k_case_box_242(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_245(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_248(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_251(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_254(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_257(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_958(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [8:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [8:0] z;
  wire [6:0] ctl;
  wire [8:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [8:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[8]), .sel1 (ctl[5]), .data1
       (in_1[8]), .sel2 (ctl[4]), .data2 (in_2[8]), .sel3 (ctl[3]),
       .data3 (in_3[8]), .sel4 (ctl[2]), .data4 (in_4[8]), .sel5
       (ctl[1]), .data5 (in_5[8]), .sel6 (ctl[0]), .data6 (in_6[8]), .z
       (z[8]));
  CDN_mux7 g10(.sel0 (ctl[6]), .data0 (in_0[7]), .sel1 (ctl[5]), .data1
       (in_1[7]), .sel2 (ctl[4]), .data2 (in_2[7]), .sel3 (ctl[3]),
       .data3 (in_3[7]), .sel4 (ctl[2]), .data4 (in_4[7]), .sel5
       (ctl[1]), .data5 (in_5[7]), .sel6 (ctl[0]), .data6 (in_6[7]), .z
       (z[7]));
  CDN_mux7 g11(.sel0 (ctl[6]), .data0 (in_0[6]), .sel1 (ctl[5]), .data1
       (in_1[6]), .sel2 (ctl[4]), .data2 (in_2[6]), .sel3 (ctl[3]),
       .data3 (in_3[6]), .sel4 (ctl[2]), .data4 (in_4[6]), .sel5
       (ctl[1]), .data5 (in_5[6]), .sel6 (ctl[0]), .data6 (in_6[6]), .z
       (z[6]));
  CDN_mux7 g12(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g13(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g14(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g15(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g16(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g17(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_case_box_260(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_976(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [5:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [5:0] z;
  wire [7:0] ctl;
  wire [5:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [5:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[5]), .sel1 (ctl[6]), .data1
       (in_1[5]), .sel2 (ctl[5]), .data2 (in_2[5]), .sel3 (ctl[4]),
       .data3 (in_3[5]), .sel4 (ctl[3]), .data4 (in_4[5]), .sel5
       (ctl[2]), .data5 (in_5[5]), .sel6 (ctl[1]), .data6 (in_6[5]),
       .sel7 (ctl[0]), .data7 (in_7[5]), .z (z[5]));
  CDN_mux8 g7(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g8(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g9(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g10(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g11(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_bmux_981(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [2:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [2:0] z;
  wire [2:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [2:0] z;
  CDN_bmux8 g1(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .z (z[2]));
  CDN_bmux8 g2(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .z (z[1]));
  CDN_bmux8 g3(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_266(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_269(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_992(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input [10:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  output [10:0] z;
  wire [11:0] ctl;
  wire [10:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  wire [10:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[10]), .sel1 (ctl[10]),
       .data1 (in_1[10]), .sel2 (ctl[9]), .data2 (in_2[10]), .sel3
       (ctl[8]), .data3 (in_3[10]), .sel4 (ctl[7]), .data4 (in_4[10]),
       .sel5 (ctl[6]), .data5 (in_5[10]), .sel6 (ctl[5]), .data6
       (in_6[10]), .sel7 (ctl[4]), .data7 (in_7[10]), .sel8 (ctl[3]),
       .data8 (in_8[10]), .sel9 (ctl[2]), .data9 (in_9[10]), .sel10
       (ctl[1]), .data10 (in_10[10]), .sel11 (ctl[0]), .data11
       (in_11[10]), .z (z[10]));
  CDN_mux12 g12(.sel0 (ctl[11]), .data0 (in_0[9]), .sel1 (ctl[10]),
       .data1 (in_1[9]), .sel2 (ctl[9]), .data2 (in_2[9]), .sel3
       (ctl[8]), .data3 (in_3[9]), .sel4 (ctl[7]), .data4 (in_4[9]),
       .sel5 (ctl[6]), .data5 (in_5[9]), .sel6 (ctl[5]), .data6
       (in_6[9]), .sel7 (ctl[4]), .data7 (in_7[9]), .sel8 (ctl[3]),
       .data8 (in_8[9]), .sel9 (ctl[2]), .data9 (in_9[9]), .sel10
       (ctl[1]), .data10 (in_10[9]), .sel11 (ctl[0]), .data11
       (in_11[9]), .z (z[9]));
  CDN_mux12 g13(.sel0 (ctl[11]), .data0 (in_0[8]), .sel1 (ctl[10]),
       .data1 (in_1[8]), .sel2 (ctl[9]), .data2 (in_2[8]), .sel3
       (ctl[8]), .data3 (in_3[8]), .sel4 (ctl[7]), .data4 (in_4[8]),
       .sel5 (ctl[6]), .data5 (in_5[8]), .sel6 (ctl[5]), .data6
       (in_6[8]), .sel7 (ctl[4]), .data7 (in_7[8]), .sel8 (ctl[3]),
       .data8 (in_8[8]), .sel9 (ctl[2]), .data9 (in_9[8]), .sel10
       (ctl[1]), .data10 (in_10[8]), .sel11 (ctl[0]), .data11
       (in_11[8]), .z (z[8]));
  CDN_mux12 g14(.sel0 (ctl[11]), .data0 (in_0[7]), .sel1 (ctl[10]),
       .data1 (in_1[7]), .sel2 (ctl[9]), .data2 (in_2[7]), .sel3
       (ctl[8]), .data3 (in_3[7]), .sel4 (ctl[7]), .data4 (in_4[7]),
       .sel5 (ctl[6]), .data5 (in_5[7]), .sel6 (ctl[5]), .data6
       (in_6[7]), .sel7 (ctl[4]), .data7 (in_7[7]), .sel8 (ctl[3]),
       .data8 (in_8[7]), .sel9 (ctl[2]), .data9 (in_9[7]), .sel10
       (ctl[1]), .data10 (in_10[7]), .sel11 (ctl[0]), .data11
       (in_11[7]), .z (z[7]));
  CDN_mux12 g15(.sel0 (ctl[11]), .data0 (in_0[6]), .sel1 (ctl[10]),
       .data1 (in_1[6]), .sel2 (ctl[9]), .data2 (in_2[6]), .sel3
       (ctl[8]), .data3 (in_3[6]), .sel4 (ctl[7]), .data4 (in_4[6]),
       .sel5 (ctl[6]), .data5 (in_5[6]), .sel6 (ctl[5]), .data6
       (in_6[6]), .sel7 (ctl[4]), .data7 (in_7[6]), .sel8 (ctl[3]),
       .data8 (in_8[6]), .sel9 (ctl[2]), .data9 (in_9[6]), .sel10
       (ctl[1]), .data10 (in_10[6]), .sel11 (ctl[0]), .data11
       (in_11[6]), .z (z[6]));
  CDN_mux12 g16(.sel0 (ctl[11]), .data0 (in_0[5]), .sel1 (ctl[10]),
       .data1 (in_1[5]), .sel2 (ctl[9]), .data2 (in_2[5]), .sel3
       (ctl[8]), .data3 (in_3[5]), .sel4 (ctl[7]), .data4 (in_4[5]),
       .sel5 (ctl[6]), .data5 (in_5[5]), .sel6 (ctl[5]), .data6
       (in_6[5]), .sel7 (ctl[4]), .data7 (in_7[5]), .sel8 (ctl[3]),
       .data8 (in_8[5]), .sel9 (ctl[2]), .data9 (in_9[5]), .sel10
       (ctl[1]), .data10 (in_10[5]), .sel11 (ctl[0]), .data11
       (in_11[5]), .z (z[5]));
  CDN_mux12 g17(.sel0 (ctl[11]), .data0 (in_0[4]), .sel1 (ctl[10]),
       .data1 (in_1[4]), .sel2 (ctl[9]), .data2 (in_2[4]), .sel3
       (ctl[8]), .data3 (in_3[4]), .sel4 (ctl[7]), .data4 (in_4[4]),
       .sel5 (ctl[6]), .data5 (in_5[4]), .sel6 (ctl[5]), .data6
       (in_6[4]), .sel7 (ctl[4]), .data7 (in_7[4]), .sel8 (ctl[3]),
       .data8 (in_8[4]), .sel9 (ctl[2]), .data9 (in_9[4]), .sel10
       (ctl[1]), .data10 (in_10[4]), .sel11 (ctl[0]), .data11
       (in_11[4]), .z (z[4]));
  CDN_mux12 g18(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g19(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g20(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g21(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_case_box_272(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_1002(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7,
       in_8, in_9, in_10, in_11;
  output [11:0] z;
  wire [11:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7,
       in_8, in_9, in_10, in_11;
  wire [11:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[11]), .sel1 (ctl[10]),
       .data1 (in_1[11]), .sel2 (ctl[9]), .data2 (in_2[11]), .sel3
       (ctl[8]), .data3 (in_3[11]), .sel4 (ctl[7]), .data4 (in_4[11]),
       .sel5 (ctl[6]), .data5 (in_5[11]), .sel6 (ctl[5]), .data6
       (in_6[11]), .sel7 (ctl[4]), .data7 (in_7[11]), .sel8 (ctl[3]),
       .data8 (in_8[11]), .sel9 (ctl[2]), .data9 (in_9[11]), .sel10
       (ctl[1]), .data10 (in_10[11]), .sel11 (ctl[0]), .data11
       (in_11[11]), .z (z[11]));
  CDN_mux12 g13(.sel0 (ctl[11]), .data0 (in_0[10]), .sel1 (ctl[10]),
       .data1 (in_1[10]), .sel2 (ctl[9]), .data2 (in_2[10]), .sel3
       (ctl[8]), .data3 (in_3[10]), .sel4 (ctl[7]), .data4 (in_4[10]),
       .sel5 (ctl[6]), .data5 (in_5[10]), .sel6 (ctl[5]), .data6
       (in_6[10]), .sel7 (ctl[4]), .data7 (in_7[10]), .sel8 (ctl[3]),
       .data8 (in_8[10]), .sel9 (ctl[2]), .data9 (in_9[10]), .sel10
       (ctl[1]), .data10 (in_10[10]), .sel11 (ctl[0]), .data11
       (in_11[10]), .z (z[10]));
  CDN_mux12 g14(.sel0 (ctl[11]), .data0 (in_0[9]), .sel1 (ctl[10]),
       .data1 (in_1[9]), .sel2 (ctl[9]), .data2 (in_2[9]), .sel3
       (ctl[8]), .data3 (in_3[9]), .sel4 (ctl[7]), .data4 (in_4[9]),
       .sel5 (ctl[6]), .data5 (in_5[9]), .sel6 (ctl[5]), .data6
       (in_6[9]), .sel7 (ctl[4]), .data7 (in_7[9]), .sel8 (ctl[3]),
       .data8 (in_8[9]), .sel9 (ctl[2]), .data9 (in_9[9]), .sel10
       (ctl[1]), .data10 (in_10[9]), .sel11 (ctl[0]), .data11
       (in_11[9]), .z (z[9]));
  CDN_mux12 g15(.sel0 (ctl[11]), .data0 (in_0[8]), .sel1 (ctl[10]),
       .data1 (in_1[8]), .sel2 (ctl[9]), .data2 (in_2[8]), .sel3
       (ctl[8]), .data3 (in_3[8]), .sel4 (ctl[7]), .data4 (in_4[8]),
       .sel5 (ctl[6]), .data5 (in_5[8]), .sel6 (ctl[5]), .data6
       (in_6[8]), .sel7 (ctl[4]), .data7 (in_7[8]), .sel8 (ctl[3]),
       .data8 (in_8[8]), .sel9 (ctl[2]), .data9 (in_9[8]), .sel10
       (ctl[1]), .data10 (in_10[8]), .sel11 (ctl[0]), .data11
       (in_11[8]), .z (z[8]));
  CDN_mux12 g16(.sel0 (ctl[11]), .data0 (in_0[7]), .sel1 (ctl[10]),
       .data1 (in_1[7]), .sel2 (ctl[9]), .data2 (in_2[7]), .sel3
       (ctl[8]), .data3 (in_3[7]), .sel4 (ctl[7]), .data4 (in_4[7]),
       .sel5 (ctl[6]), .data5 (in_5[7]), .sel6 (ctl[5]), .data6
       (in_6[7]), .sel7 (ctl[4]), .data7 (in_7[7]), .sel8 (ctl[3]),
       .data8 (in_8[7]), .sel9 (ctl[2]), .data9 (in_9[7]), .sel10
       (ctl[1]), .data10 (in_10[7]), .sel11 (ctl[0]), .data11
       (in_11[7]), .z (z[7]));
  CDN_mux12 g17(.sel0 (ctl[11]), .data0 (in_0[6]), .sel1 (ctl[10]),
       .data1 (in_1[6]), .sel2 (ctl[9]), .data2 (in_2[6]), .sel3
       (ctl[8]), .data3 (in_3[6]), .sel4 (ctl[7]), .data4 (in_4[6]),
       .sel5 (ctl[6]), .data5 (in_5[6]), .sel6 (ctl[5]), .data6
       (in_6[6]), .sel7 (ctl[4]), .data7 (in_7[6]), .sel8 (ctl[3]),
       .data8 (in_8[6]), .sel9 (ctl[2]), .data9 (in_9[6]), .sel10
       (ctl[1]), .data10 (in_10[6]), .sel11 (ctl[0]), .data11
       (in_11[6]), .z (z[6]));
  CDN_mux12 g18(.sel0 (ctl[11]), .data0 (in_0[5]), .sel1 (ctl[10]),
       .data1 (in_1[5]), .sel2 (ctl[9]), .data2 (in_2[5]), .sel3
       (ctl[8]), .data3 (in_3[5]), .sel4 (ctl[7]), .data4 (in_4[5]),
       .sel5 (ctl[6]), .data5 (in_5[5]), .sel6 (ctl[5]), .data6
       (in_6[5]), .sel7 (ctl[4]), .data7 (in_7[5]), .sel8 (ctl[3]),
       .data8 (in_8[5]), .sel9 (ctl[2]), .data9 (in_9[5]), .sel10
       (ctl[1]), .data10 (in_10[5]), .sel11 (ctl[0]), .data11
       (in_11[5]), .z (z[5]));
  CDN_mux12 g19(.sel0 (ctl[11]), .data0 (in_0[4]), .sel1 (ctl[10]),
       .data1 (in_1[4]), .sel2 (ctl[9]), .data2 (in_2[4]), .sel3
       (ctl[8]), .data3 (in_3[4]), .sel4 (ctl[7]), .data4 (in_4[4]),
       .sel5 (ctl[6]), .data5 (in_5[4]), .sel6 (ctl[5]), .data6
       (in_6[4]), .sel7 (ctl[4]), .data7 (in_7[4]), .sel8 (ctl[3]),
       .data8 (in_8[4]), .sel9 (ctl[2]), .data9 (in_9[4]), .sel10
       (ctl[1]), .data10 (in_10[4]), .sel11 (ctl[0]), .data11
       (in_11[4]), .z (z[4]));
  CDN_mux12 g20(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g21(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g22(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g23(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_case_box_275(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_278(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_281(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_284(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_287(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_1062(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [3:0] z;
  wire [7:0] ctl;
  wire [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [3:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g5(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g6(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g7(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_293(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_296(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_299(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_302(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_305(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_308(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_311(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_314(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_320(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_323(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_326(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_329(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_332(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_335(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_338(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_341(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_1224(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [4:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [4:0] z;
  wire [7:0] ctl;
  wire [4:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [4:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g6(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g7(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g8(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g9(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_bmux_1228(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [2:0] ctl;
  input [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [3:0] z;
  wire [2:0] ctl;
  wire [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [3:0] z;
  CDN_bmux8 g1(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .z (z[3]));
  CDN_bmux8 g2(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .z (z[2]));
  CDN_bmux8 g3(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .z (z[1]));
  CDN_bmux8 g4(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_347(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_350(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_353(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_356(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_359(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_362(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_365(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_368(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_bmux_1313(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, z);
  input [3:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15;
  output [9:0] z;
  wire [3:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15;
  wire [9:0] z;
  CDN_bmux16 g1(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .sel2
       (ctl[2]), .data4 (in_4[9]), .data5 (in_5[9]), .data6 (in_6[9]),
       .data7 (in_7[9]), .sel3 (ctl[3]), .data8 (in_8[9]), .data9
       (in_9[9]), .data10 (in_10[9]), .data11 (in_11[9]), .data12
       (in_12[9]), .data13 (in_13[9]), .data14 (in_14[9]), .data15
       (in_15[9]), .z (z[9]));
  CDN_bmux16 g2(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .sel2
       (ctl[2]), .data4 (in_4[8]), .data5 (in_5[8]), .data6 (in_6[8]),
       .data7 (in_7[8]), .sel3 (ctl[3]), .data8 (in_8[8]), .data9
       (in_9[8]), .data10 (in_10[8]), .data11 (in_11[8]), .data12
       (in_12[8]), .data13 (in_13[8]), .data14 (in_14[8]), .data15
       (in_15[8]), .z (z[8]));
  CDN_bmux16 g3(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .data7 (in_7[7]), .sel3 (ctl[3]), .data8 (in_8[7]), .data9
       (in_9[7]), .data10 (in_10[7]), .data11 (in_11[7]), .data12
       (in_12[7]), .data13 (in_13[7]), .data14 (in_14[7]), .data15
       (in_15[7]), .z (z[7]));
  CDN_bmux16 g4(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .data7 (in_7[6]), .sel3 (ctl[3]), .data8 (in_8[6]), .data9
       (in_9[6]), .data10 (in_10[6]), .data11 (in_11[6]), .data12
       (in_12[6]), .data13 (in_13[6]), .data14 (in_14[6]), .data15
       (in_15[6]), .z (z[6]));
  CDN_bmux16 g5(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .data7 (in_7[5]), .sel3 (ctl[3]), .data8 (in_8[5]), .data9
       (in_9[5]), .data10 (in_10[5]), .data11 (in_11[5]), .data12
       (in_12[5]), .data13 (in_13[5]), .data14 (in_14[5]), .data15
       (in_15[5]), .z (z[5]));
  CDN_bmux16 g6(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .data7 (in_7[4]), .sel3 (ctl[3]), .data8 (in_8[4]), .data9
       (in_9[4]), .data10 (in_10[4]), .data11 (in_11[4]), .data12
       (in_12[4]), .data13 (in_13[4]), .data14 (in_14[4]), .data15
       (in_15[4]), .z (z[4]));
  CDN_bmux16 g7(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .sel3 (ctl[3]), .data8 (in_8[3]), .data9
       (in_9[3]), .data10 (in_10[3]), .data11 (in_11[3]), .data12
       (in_12[3]), .data13 (in_13[3]), .data14 (in_14[3]), .data15
       (in_15[3]), .z (z[3]));
  CDN_bmux16 g8(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .sel3 (ctl[3]), .data8 (in_8[2]), .data9
       (in_9[2]), .data10 (in_10[2]), .data11 (in_11[2]), .data12
       (in_12[2]), .data13 (in_13[2]), .data14 (in_14[2]), .data15
       (in_15[2]), .z (z[2]));
  CDN_bmux16 g9(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .sel3 (ctl[3]), .data8 (in_8[1]), .data9
       (in_9[1]), .data10 (in_10[1]), .data11 (in_11[1]), .data12
       (in_12[1]), .data13 (in_13[1]), .data14 (in_14[1]), .data15
       (in_15[1]), .z (z[1]));
  CDN_bmux16 g10(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .sel3 (ctl[3]), .data8 (in_8[0]), .data9
       (in_9[0]), .data10 (in_10[0]), .data11 (in_11[0]), .data12
       (in_12[0]), .data13 (in_13[0]), .data14 (in_14[0]), .data15
       (in_15[0]), .z (z[0]));
endmodule

module fx68k_mux_1316(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [4:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [4:0] z;
  wire [6:0] ctl;
  wire [4:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [4:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g6(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g7(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g8(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g9(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_bmux_1352(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, z);
  input [3:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  output [9:0] z;
  wire [3:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  wire [9:0] z;
  CDN_bmux9 g1(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .sel2
       (ctl[2]), .data4 (in_4[9]), .data5 (in_5[9]), .data6 (in_6[9]),
       .data7 (in_7[9]), .sel3 (ctl[3]), .data8 (in_8[9]), .z (z[9]));
  CDN_bmux9 g2(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .sel2
       (ctl[2]), .data4 (in_4[8]), .data5 (in_5[8]), .data6 (in_6[8]),
       .data7 (in_7[8]), .sel3 (ctl[3]), .data8 (in_8[8]), .z (z[8]));
  CDN_bmux9 g3(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .data7 (in_7[7]), .sel3 (ctl[3]), .data8 (in_8[7]), .z (z[7]));
  CDN_bmux9 g4(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .data7 (in_7[6]), .sel3 (ctl[3]), .data8 (in_8[6]), .z (z[6]));
  CDN_bmux9 g5(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .data7 (in_7[5]), .sel3 (ctl[3]), .data8 (in_8[5]), .z (z[5]));
  CDN_bmux9 g6(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .data7 (in_7[4]), .sel3 (ctl[3]), .data8 (in_8[4]), .z (z[4]));
  CDN_bmux9 g7(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .sel3 (ctl[3]), .data8 (in_8[3]), .z (z[3]));
  CDN_bmux9 g8(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .sel3 (ctl[3]), .data8 (in_8[2]), .z (z[2]));
  CDN_bmux9 g9(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .sel3 (ctl[3]), .data8 (in_8[1]), .z (z[1]));
  CDN_bmux9 g10(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .sel3 (ctl[3]), .data8 (in_8[0]), .z (z[0]));
endmodule

module fx68k_case_box_374(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_1354(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input [17:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [17:0] z;
  wire [7:0] ctl;
  wire [17:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [17:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[17]), .sel1 (ctl[6]), .data1
       (in_1[17]), .sel2 (ctl[5]), .data2 (in_2[17]), .sel3 (ctl[4]),
       .data3 (in_3[17]), .sel4 (ctl[3]), .data4 (in_4[17]), .sel5
       (ctl[2]), .data5 (in_5[17]), .sel6 (ctl[1]), .data6 (in_6[17]),
       .sel7 (ctl[0]), .data7 (in_7[17]), .z (z[17]));
  CDN_mux8 g19(.sel0 (ctl[7]), .data0 (in_0[16]), .sel1 (ctl[6]),
       .data1 (in_1[16]), .sel2 (ctl[5]), .data2 (in_2[16]), .sel3
       (ctl[4]), .data3 (in_3[16]), .sel4 (ctl[3]), .data4 (in_4[16]),
       .sel5 (ctl[2]), .data5 (in_5[16]), .sel6 (ctl[1]), .data6
       (in_6[16]), .sel7 (ctl[0]), .data7 (in_7[16]), .z (z[16]));
  CDN_mux8 g20(.sel0 (ctl[7]), .data0 (in_0[15]), .sel1 (ctl[6]),
       .data1 (in_1[15]), .sel2 (ctl[5]), .data2 (in_2[15]), .sel3
       (ctl[4]), .data3 (in_3[15]), .sel4 (ctl[3]), .data4 (in_4[15]),
       .sel5 (ctl[2]), .data5 (in_5[15]), .sel6 (ctl[1]), .data6
       (in_6[15]), .sel7 (ctl[0]), .data7 (in_7[15]), .z (z[15]));
  CDN_mux8 g21(.sel0 (ctl[7]), .data0 (in_0[14]), .sel1 (ctl[6]),
       .data1 (in_1[14]), .sel2 (ctl[5]), .data2 (in_2[14]), .sel3
       (ctl[4]), .data3 (in_3[14]), .sel4 (ctl[3]), .data4 (in_4[14]),
       .sel5 (ctl[2]), .data5 (in_5[14]), .sel6 (ctl[1]), .data6
       (in_6[14]), .sel7 (ctl[0]), .data7 (in_7[14]), .z (z[14]));
  CDN_mux8 g22(.sel0 (ctl[7]), .data0 (in_0[13]), .sel1 (ctl[6]),
       .data1 (in_1[13]), .sel2 (ctl[5]), .data2 (in_2[13]), .sel3
       (ctl[4]), .data3 (in_3[13]), .sel4 (ctl[3]), .data4 (in_4[13]),
       .sel5 (ctl[2]), .data5 (in_5[13]), .sel6 (ctl[1]), .data6
       (in_6[13]), .sel7 (ctl[0]), .data7 (in_7[13]), .z (z[13]));
  CDN_mux8 g23(.sel0 (ctl[7]), .data0 (in_0[12]), .sel1 (ctl[6]),
       .data1 (in_1[12]), .sel2 (ctl[5]), .data2 (in_2[12]), .sel3
       (ctl[4]), .data3 (in_3[12]), .sel4 (ctl[3]), .data4 (in_4[12]),
       .sel5 (ctl[2]), .data5 (in_5[12]), .sel6 (ctl[1]), .data6
       (in_6[12]), .sel7 (ctl[0]), .data7 (in_7[12]), .z (z[12]));
  CDN_mux8 g24(.sel0 (ctl[7]), .data0 (in_0[11]), .sel1 (ctl[6]),
       .data1 (in_1[11]), .sel2 (ctl[5]), .data2 (in_2[11]), .sel3
       (ctl[4]), .data3 (in_3[11]), .sel4 (ctl[3]), .data4 (in_4[11]),
       .sel5 (ctl[2]), .data5 (in_5[11]), .sel6 (ctl[1]), .data6
       (in_6[11]), .sel7 (ctl[0]), .data7 (in_7[11]), .z (z[11]));
  CDN_mux8 g25(.sel0 (ctl[7]), .data0 (in_0[10]), .sel1 (ctl[6]),
       .data1 (in_1[10]), .sel2 (ctl[5]), .data2 (in_2[10]), .sel3
       (ctl[4]), .data3 (in_3[10]), .sel4 (ctl[3]), .data4 (in_4[10]),
       .sel5 (ctl[2]), .data5 (in_5[10]), .sel6 (ctl[1]), .data6
       (in_6[10]), .sel7 (ctl[0]), .data7 (in_7[10]), .z (z[10]));
  CDN_mux8 g26(.sel0 (ctl[7]), .data0 (in_0[9]), .sel1 (ctl[6]), .data1
       (in_1[9]), .sel2 (ctl[5]), .data2 (in_2[9]), .sel3 (ctl[4]),
       .data3 (in_3[9]), .sel4 (ctl[3]), .data4 (in_4[9]), .sel5
       (ctl[2]), .data5 (in_5[9]), .sel6 (ctl[1]), .data6 (in_6[9]),
       .sel7 (ctl[0]), .data7 (in_7[9]), .z (z[9]));
  CDN_mux8 g27(.sel0 (ctl[7]), .data0 (in_0[8]), .sel1 (ctl[6]), .data1
       (in_1[8]), .sel2 (ctl[5]), .data2 (in_2[8]), .sel3 (ctl[4]),
       .data3 (in_3[8]), .sel4 (ctl[3]), .data4 (in_4[8]), .sel5
       (ctl[2]), .data5 (in_5[8]), .sel6 (ctl[1]), .data6 (in_6[8]),
       .sel7 (ctl[0]), .data7 (in_7[8]), .z (z[8]));
  CDN_mux8 g28(.sel0 (ctl[7]), .data0 (in_0[7]), .sel1 (ctl[6]), .data1
       (in_1[7]), .sel2 (ctl[5]), .data2 (in_2[7]), .sel3 (ctl[4]),
       .data3 (in_3[7]), .sel4 (ctl[3]), .data4 (in_4[7]), .sel5
       (ctl[2]), .data5 (in_5[7]), .sel6 (ctl[1]), .data6 (in_6[7]),
       .sel7 (ctl[0]), .data7 (in_7[7]), .z (z[7]));
  CDN_mux8 g29(.sel0 (ctl[7]), .data0 (in_0[6]), .sel1 (ctl[6]), .data1
       (in_1[6]), .sel2 (ctl[5]), .data2 (in_2[6]), .sel3 (ctl[4]),
       .data3 (in_3[6]), .sel4 (ctl[3]), .data4 (in_4[6]), .sel5
       (ctl[2]), .data5 (in_5[6]), .sel6 (ctl[1]), .data6 (in_6[6]),
       .sel7 (ctl[0]), .data7 (in_7[6]), .z (z[6]));
  CDN_mux8 g30(.sel0 (ctl[7]), .data0 (in_0[5]), .sel1 (ctl[6]), .data1
       (in_1[5]), .sel2 (ctl[5]), .data2 (in_2[5]), .sel3 (ctl[4]),
       .data3 (in_3[5]), .sel4 (ctl[3]), .data4 (in_4[5]), .sel5
       (ctl[2]), .data5 (in_5[5]), .sel6 (ctl[1]), .data6 (in_6[5]),
       .sel7 (ctl[0]), .data7 (in_7[5]), .z (z[5]));
  CDN_mux8 g31(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g32(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g33(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g34(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g35(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_case_box_377(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_1371(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [17:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [17:0] z;
  wire [6:0] ctl;
  wire [17:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [17:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[17]), .sel1 (ctl[5]), .data1
       (in_1[17]), .sel2 (ctl[4]), .data2 (in_2[17]), .sel3 (ctl[3]),
       .data3 (in_3[17]), .sel4 (ctl[2]), .data4 (in_4[17]), .sel5
       (ctl[1]), .data5 (in_5[17]), .sel6 (ctl[0]), .data6 (in_6[17]),
       .z (z[17]));
  CDN_mux7 g19(.sel0 (ctl[6]), .data0 (in_0[16]), .sel1 (ctl[5]),
       .data1 (in_1[16]), .sel2 (ctl[4]), .data2 (in_2[16]), .sel3
       (ctl[3]), .data3 (in_3[16]), .sel4 (ctl[2]), .data4 (in_4[16]),
       .sel5 (ctl[1]), .data5 (in_5[16]), .sel6 (ctl[0]), .data6
       (in_6[16]), .z (z[16]));
  CDN_mux7 g20(.sel0 (ctl[6]), .data0 (in_0[15]), .sel1 (ctl[5]),
       .data1 (in_1[15]), .sel2 (ctl[4]), .data2 (in_2[15]), .sel3
       (ctl[3]), .data3 (in_3[15]), .sel4 (ctl[2]), .data4 (in_4[15]),
       .sel5 (ctl[1]), .data5 (in_5[15]), .sel6 (ctl[0]), .data6
       (in_6[15]), .z (z[15]));
  CDN_mux7 g21(.sel0 (ctl[6]), .data0 (in_0[14]), .sel1 (ctl[5]),
       .data1 (in_1[14]), .sel2 (ctl[4]), .data2 (in_2[14]), .sel3
       (ctl[3]), .data3 (in_3[14]), .sel4 (ctl[2]), .data4 (in_4[14]),
       .sel5 (ctl[1]), .data5 (in_5[14]), .sel6 (ctl[0]), .data6
       (in_6[14]), .z (z[14]));
  CDN_mux7 g22(.sel0 (ctl[6]), .data0 (in_0[13]), .sel1 (ctl[5]),
       .data1 (in_1[13]), .sel2 (ctl[4]), .data2 (in_2[13]), .sel3
       (ctl[3]), .data3 (in_3[13]), .sel4 (ctl[2]), .data4 (in_4[13]),
       .sel5 (ctl[1]), .data5 (in_5[13]), .sel6 (ctl[0]), .data6
       (in_6[13]), .z (z[13]));
  CDN_mux7 g23(.sel0 (ctl[6]), .data0 (in_0[12]), .sel1 (ctl[5]),
       .data1 (in_1[12]), .sel2 (ctl[4]), .data2 (in_2[12]), .sel3
       (ctl[3]), .data3 (in_3[12]), .sel4 (ctl[2]), .data4 (in_4[12]),
       .sel5 (ctl[1]), .data5 (in_5[12]), .sel6 (ctl[0]), .data6
       (in_6[12]), .z (z[12]));
  CDN_mux7 g24(.sel0 (ctl[6]), .data0 (in_0[11]), .sel1 (ctl[5]),
       .data1 (in_1[11]), .sel2 (ctl[4]), .data2 (in_2[11]), .sel3
       (ctl[3]), .data3 (in_3[11]), .sel4 (ctl[2]), .data4 (in_4[11]),
       .sel5 (ctl[1]), .data5 (in_5[11]), .sel6 (ctl[0]), .data6
       (in_6[11]), .z (z[11]));
  CDN_mux7 g25(.sel0 (ctl[6]), .data0 (in_0[10]), .sel1 (ctl[5]),
       .data1 (in_1[10]), .sel2 (ctl[4]), .data2 (in_2[10]), .sel3
       (ctl[3]), .data3 (in_3[10]), .sel4 (ctl[2]), .data4 (in_4[10]),
       .sel5 (ctl[1]), .data5 (in_5[10]), .sel6 (ctl[0]), .data6
       (in_6[10]), .z (z[10]));
  CDN_mux7 g26(.sel0 (ctl[6]), .data0 (in_0[9]), .sel1 (ctl[5]), .data1
       (in_1[9]), .sel2 (ctl[4]), .data2 (in_2[9]), .sel3 (ctl[3]),
       .data3 (in_3[9]), .sel4 (ctl[2]), .data4 (in_4[9]), .sel5
       (ctl[1]), .data5 (in_5[9]), .sel6 (ctl[0]), .data6 (in_6[9]), .z
       (z[9]));
  CDN_mux7 g27(.sel0 (ctl[6]), .data0 (in_0[8]), .sel1 (ctl[5]), .data1
       (in_1[8]), .sel2 (ctl[4]), .data2 (in_2[8]), .sel3 (ctl[3]),
       .data3 (in_3[8]), .sel4 (ctl[2]), .data4 (in_4[8]), .sel5
       (ctl[1]), .data5 (in_5[8]), .sel6 (ctl[0]), .data6 (in_6[8]), .z
       (z[8]));
  CDN_mux7 g28(.sel0 (ctl[6]), .data0 (in_0[7]), .sel1 (ctl[5]), .data1
       (in_1[7]), .sel2 (ctl[4]), .data2 (in_2[7]), .sel3 (ctl[3]),
       .data3 (in_3[7]), .sel4 (ctl[2]), .data4 (in_4[7]), .sel5
       (ctl[1]), .data5 (in_5[7]), .sel6 (ctl[0]), .data6 (in_6[7]), .z
       (z[7]));
  CDN_mux7 g29(.sel0 (ctl[6]), .data0 (in_0[6]), .sel1 (ctl[5]), .data1
       (in_1[6]), .sel2 (ctl[4]), .data2 (in_2[6]), .sel3 (ctl[3]),
       .data3 (in_3[6]), .sel4 (ctl[2]), .data4 (in_4[6]), .sel5
       (ctl[1]), .data5 (in_5[6]), .sel6 (ctl[0]), .data6 (in_6[6]), .z
       (z[6]));
  CDN_mux7 g30(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g31(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g32(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g33(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g34(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g35(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_case_box_380(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_1388(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [18:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [18:0] z;
  wire [6:0] ctl;
  wire [18:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [18:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[18]), .sel1 (ctl[5]), .data1
       (in_1[18]), .sel2 (ctl[4]), .data2 (in_2[18]), .sel3 (ctl[3]),
       .data3 (in_3[18]), .sel4 (ctl[2]), .data4 (in_4[18]), .sel5
       (ctl[1]), .data5 (in_5[18]), .sel6 (ctl[0]), .data6 (in_6[18]),
       .z (z[18]));
  CDN_mux7 g20(.sel0 (ctl[6]), .data0 (in_0[17]), .sel1 (ctl[5]),
       .data1 (in_1[17]), .sel2 (ctl[4]), .data2 (in_2[17]), .sel3
       (ctl[3]), .data3 (in_3[17]), .sel4 (ctl[2]), .data4 (in_4[17]),
       .sel5 (ctl[1]), .data5 (in_5[17]), .sel6 (ctl[0]), .data6
       (in_6[17]), .z (z[17]));
  CDN_mux7 g21(.sel0 (ctl[6]), .data0 (in_0[16]), .sel1 (ctl[5]),
       .data1 (in_1[16]), .sel2 (ctl[4]), .data2 (in_2[16]), .sel3
       (ctl[3]), .data3 (in_3[16]), .sel4 (ctl[2]), .data4 (in_4[16]),
       .sel5 (ctl[1]), .data5 (in_5[16]), .sel6 (ctl[0]), .data6
       (in_6[16]), .z (z[16]));
  CDN_mux7 g22(.sel0 (ctl[6]), .data0 (in_0[15]), .sel1 (ctl[5]),
       .data1 (in_1[15]), .sel2 (ctl[4]), .data2 (in_2[15]), .sel3
       (ctl[3]), .data3 (in_3[15]), .sel4 (ctl[2]), .data4 (in_4[15]),
       .sel5 (ctl[1]), .data5 (in_5[15]), .sel6 (ctl[0]), .data6
       (in_6[15]), .z (z[15]));
  CDN_mux7 g23(.sel0 (ctl[6]), .data0 (in_0[14]), .sel1 (ctl[5]),
       .data1 (in_1[14]), .sel2 (ctl[4]), .data2 (in_2[14]), .sel3
       (ctl[3]), .data3 (in_3[14]), .sel4 (ctl[2]), .data4 (in_4[14]),
       .sel5 (ctl[1]), .data5 (in_5[14]), .sel6 (ctl[0]), .data6
       (in_6[14]), .z (z[14]));
  CDN_mux7 g24(.sel0 (ctl[6]), .data0 (in_0[13]), .sel1 (ctl[5]),
       .data1 (in_1[13]), .sel2 (ctl[4]), .data2 (in_2[13]), .sel3
       (ctl[3]), .data3 (in_3[13]), .sel4 (ctl[2]), .data4 (in_4[13]),
       .sel5 (ctl[1]), .data5 (in_5[13]), .sel6 (ctl[0]), .data6
       (in_6[13]), .z (z[13]));
  CDN_mux7 g25(.sel0 (ctl[6]), .data0 (in_0[12]), .sel1 (ctl[5]),
       .data1 (in_1[12]), .sel2 (ctl[4]), .data2 (in_2[12]), .sel3
       (ctl[3]), .data3 (in_3[12]), .sel4 (ctl[2]), .data4 (in_4[12]),
       .sel5 (ctl[1]), .data5 (in_5[12]), .sel6 (ctl[0]), .data6
       (in_6[12]), .z (z[12]));
  CDN_mux7 g26(.sel0 (ctl[6]), .data0 (in_0[11]), .sel1 (ctl[5]),
       .data1 (in_1[11]), .sel2 (ctl[4]), .data2 (in_2[11]), .sel3
       (ctl[3]), .data3 (in_3[11]), .sel4 (ctl[2]), .data4 (in_4[11]),
       .sel5 (ctl[1]), .data5 (in_5[11]), .sel6 (ctl[0]), .data6
       (in_6[11]), .z (z[11]));
  CDN_mux7 g27(.sel0 (ctl[6]), .data0 (in_0[10]), .sel1 (ctl[5]),
       .data1 (in_1[10]), .sel2 (ctl[4]), .data2 (in_2[10]), .sel3
       (ctl[3]), .data3 (in_3[10]), .sel4 (ctl[2]), .data4 (in_4[10]),
       .sel5 (ctl[1]), .data5 (in_5[10]), .sel6 (ctl[0]), .data6
       (in_6[10]), .z (z[10]));
  CDN_mux7 g28(.sel0 (ctl[6]), .data0 (in_0[9]), .sel1 (ctl[5]), .data1
       (in_1[9]), .sel2 (ctl[4]), .data2 (in_2[9]), .sel3 (ctl[3]),
       .data3 (in_3[9]), .sel4 (ctl[2]), .data4 (in_4[9]), .sel5
       (ctl[1]), .data5 (in_5[9]), .sel6 (ctl[0]), .data6 (in_6[9]), .z
       (z[9]));
  CDN_mux7 g29(.sel0 (ctl[6]), .data0 (in_0[8]), .sel1 (ctl[5]), .data1
       (in_1[8]), .sel2 (ctl[4]), .data2 (in_2[8]), .sel3 (ctl[3]),
       .data3 (in_3[8]), .sel4 (ctl[2]), .data4 (in_4[8]), .sel5
       (ctl[1]), .data5 (in_5[8]), .sel6 (ctl[0]), .data6 (in_6[8]), .z
       (z[8]));
  CDN_mux7 g30(.sel0 (ctl[6]), .data0 (in_0[7]), .sel1 (ctl[5]), .data1
       (in_1[7]), .sel2 (ctl[4]), .data2 (in_2[7]), .sel3 (ctl[3]),
       .data3 (in_3[7]), .sel4 (ctl[2]), .data4 (in_4[7]), .sel5
       (ctl[1]), .data5 (in_5[7]), .sel6 (ctl[0]), .data6 (in_6[7]), .z
       (z[7]));
  CDN_mux7 g31(.sel0 (ctl[6]), .data0 (in_0[6]), .sel1 (ctl[5]), .data1
       (in_1[6]), .sel2 (ctl[4]), .data2 (in_2[6]), .sel3 (ctl[3]),
       .data3 (in_3[6]), .sel4 (ctl[2]), .data4 (in_4[6]), .sel5
       (ctl[1]), .data5 (in_5[6]), .sel6 (ctl[0]), .data6 (in_6[6]), .z
       (z[6]));
  CDN_mux7 g32(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g33(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g34(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g35(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g36(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g37(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_case_box_383(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_386(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_mux_1423(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [16:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [16:0] z;
  wire [6:0] ctl;
  wire [16:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [16:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[16]), .sel1 (ctl[5]), .data1
       (in_1[16]), .sel2 (ctl[4]), .data2 (in_2[16]), .sel3 (ctl[3]),
       .data3 (in_3[16]), .sel4 (ctl[2]), .data4 (in_4[16]), .sel5
       (ctl[1]), .data5 (in_5[16]), .sel6 (ctl[0]), .data6 (in_6[16]),
       .z (z[16]));
  CDN_mux7 g18(.sel0 (ctl[6]), .data0 (in_0[15]), .sel1 (ctl[5]),
       .data1 (in_1[15]), .sel2 (ctl[4]), .data2 (in_2[15]), .sel3
       (ctl[3]), .data3 (in_3[15]), .sel4 (ctl[2]), .data4 (in_4[15]),
       .sel5 (ctl[1]), .data5 (in_5[15]), .sel6 (ctl[0]), .data6
       (in_6[15]), .z (z[15]));
  CDN_mux7 g19(.sel0 (ctl[6]), .data0 (in_0[14]), .sel1 (ctl[5]),
       .data1 (in_1[14]), .sel2 (ctl[4]), .data2 (in_2[14]), .sel3
       (ctl[3]), .data3 (in_3[14]), .sel4 (ctl[2]), .data4 (in_4[14]),
       .sel5 (ctl[1]), .data5 (in_5[14]), .sel6 (ctl[0]), .data6
       (in_6[14]), .z (z[14]));
  CDN_mux7 g20(.sel0 (ctl[6]), .data0 (in_0[13]), .sel1 (ctl[5]),
       .data1 (in_1[13]), .sel2 (ctl[4]), .data2 (in_2[13]), .sel3
       (ctl[3]), .data3 (in_3[13]), .sel4 (ctl[2]), .data4 (in_4[13]),
       .sel5 (ctl[1]), .data5 (in_5[13]), .sel6 (ctl[0]), .data6
       (in_6[13]), .z (z[13]));
  CDN_mux7 g21(.sel0 (ctl[6]), .data0 (in_0[12]), .sel1 (ctl[5]),
       .data1 (in_1[12]), .sel2 (ctl[4]), .data2 (in_2[12]), .sel3
       (ctl[3]), .data3 (in_3[12]), .sel4 (ctl[2]), .data4 (in_4[12]),
       .sel5 (ctl[1]), .data5 (in_5[12]), .sel6 (ctl[0]), .data6
       (in_6[12]), .z (z[12]));
  CDN_mux7 g22(.sel0 (ctl[6]), .data0 (in_0[11]), .sel1 (ctl[5]),
       .data1 (in_1[11]), .sel2 (ctl[4]), .data2 (in_2[11]), .sel3
       (ctl[3]), .data3 (in_3[11]), .sel4 (ctl[2]), .data4 (in_4[11]),
       .sel5 (ctl[1]), .data5 (in_5[11]), .sel6 (ctl[0]), .data6
       (in_6[11]), .z (z[11]));
  CDN_mux7 g23(.sel0 (ctl[6]), .data0 (in_0[10]), .sel1 (ctl[5]),
       .data1 (in_1[10]), .sel2 (ctl[4]), .data2 (in_2[10]), .sel3
       (ctl[3]), .data3 (in_3[10]), .sel4 (ctl[2]), .data4 (in_4[10]),
       .sel5 (ctl[1]), .data5 (in_5[10]), .sel6 (ctl[0]), .data6
       (in_6[10]), .z (z[10]));
  CDN_mux7 g24(.sel0 (ctl[6]), .data0 (in_0[9]), .sel1 (ctl[5]), .data1
       (in_1[9]), .sel2 (ctl[4]), .data2 (in_2[9]), .sel3 (ctl[3]),
       .data3 (in_3[9]), .sel4 (ctl[2]), .data4 (in_4[9]), .sel5
       (ctl[1]), .data5 (in_5[9]), .sel6 (ctl[0]), .data6 (in_6[9]), .z
       (z[9]));
  CDN_mux7 g25(.sel0 (ctl[6]), .data0 (in_0[8]), .sel1 (ctl[5]), .data1
       (in_1[8]), .sel2 (ctl[4]), .data2 (in_2[8]), .sel3 (ctl[3]),
       .data3 (in_3[8]), .sel4 (ctl[2]), .data4 (in_4[8]), .sel5
       (ctl[1]), .data5 (in_5[8]), .sel6 (ctl[0]), .data6 (in_6[8]), .z
       (z[8]));
  CDN_mux7 g26(.sel0 (ctl[6]), .data0 (in_0[7]), .sel1 (ctl[5]), .data1
       (in_1[7]), .sel2 (ctl[4]), .data2 (in_2[7]), .sel3 (ctl[3]),
       .data3 (in_3[7]), .sel4 (ctl[2]), .data4 (in_4[7]), .sel5
       (ctl[1]), .data5 (in_5[7]), .sel6 (ctl[0]), .data6 (in_6[7]), .z
       (z[7]));
  CDN_mux7 g27(.sel0 (ctl[6]), .data0 (in_0[6]), .sel1 (ctl[5]), .data1
       (in_1[6]), .sel2 (ctl[4]), .data2 (in_2[6]), .sel3 (ctl[3]),
       .data3 (in_3[6]), .sel4 (ctl[2]), .data4 (in_4[6]), .sel5
       (ctl[1]), .data5 (in_5[6]), .sel6 (ctl[0]), .data6 (in_6[6]), .z
       (z[6]));
  CDN_mux7 g28(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g29(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g30(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g31(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g32(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g33(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_case_box_389(in_0, out_0);
  input [3:0] in_0;
  output [12:0] out_0;
  wire [3:0] in_0;
  wire [12:0] out_0;
  wire n_5, n_7, n_9, n_10, n_12, n_14, n_17, n_20;
  wire n_23, n_26, n_114, n_115;
  assign out_0[0] = 1'b0;
  nor g1 (out_0[12], n_5, n_10);
  nand g2 (n_5, n_114, n_115);
  not g3 (n_114, in_0[0]);
  not g4 (n_115, in_0[2]);
  nand g5 (n_10, n_7, n_9);
  not g6 (n_7, in_0[1]);
  not g7 (n_9, in_0[3]);
  nor g8 (out_0[11], n_10, n_12);
  nand g9 (n_12, in_0[0], n_115);
  nor g10 (out_0[10], n_5, n_14);
  nand g11 (n_14, in_0[1], n_9);
  nor g12 (out_0[9], n_12, n_14);
  nor g13 (out_0[8], in_0[0], n_17);
  nand g14 (n_17, n_7, in_0[2]);
  nor g15 (out_0[7], n_17, n_114);
  nor g16 (out_0[6], in_0[0], n_20);
  nand g17 (n_20, in_0[1], in_0[2]);
  nor g18 (out_0[5], n_20, n_114);
  nor g19 (out_0[4], in_0[0], n_23);
  nand g20 (n_23, n_7, in_0[3]);
  nor g21 (out_0[3], n_23, n_114);
  nor g22 (out_0[2], in_0[0], n_26);
  nand g23 (n_26, in_0[1], in_0[3]);
  nor g24 (out_0[1], n_26, n_114);
endmodule

module fx68k_case_box_392(in_0, out_0);
  input [2:0] in_0;
  output [7:0] out_0;
  wire [2:0] in_0;
  wire [7:0] out_0;
  wire n_6, n_8, n_9, n_11, n_14, n_54, n_55;
  nor g1 (out_0[7], n_54, n_6);
  not g2 (n_54, in_0[2]);
  nand g3 (n_6, in_0[1], n_55);
  not g4 (n_55, in_0[0]);
  nor g5 (out_0[6], in_0[2], n_9);
  nand g6 (n_9, n_8, n_55);
  not g7 (n_8, in_0[1]);
  nor g8 (out_0[5], in_0[2], n_11);
  nand g9 (n_11, n_8, in_0[0]);
  nor g10 (out_0[4], n_6, in_0[2]);
  nor g11 (out_0[3], in_0[2], n_14);
  nand g12 (n_14, in_0[1], in_0[0]);
  nor g13 (out_0[2], n_14, n_54);
  nor g14 (out_0[1], n_11, n_54);
  nor g15 (out_0[0], n_9, n_54);
endmodule

module fx68k_mux_1463(ctl, in_0, in_1, in_2, in_3, in_4, in_5, z);
  input [5:0] ctl;
  input [1:0] in_0, in_1, in_2, in_3, in_4, in_5;
  output [1:0] z;
  wire [5:0] ctl;
  wire [1:0] in_0, in_1, in_2, in_3, in_4, in_5;
  wire [1:0] z;
  CDN_mux6 g1(.sel0 (ctl[5]), .data0 (in_0[1]), .sel1 (ctl[4]), .data1
       (in_1[1]), .sel2 (ctl[3]), .data2 (in_2[1]), .sel3 (ctl[2]),
       .data3 (in_3[1]), .sel4 (ctl[1]), .data4 (in_4[1]), .sel5
       (ctl[0]), .data5 (in_5[1]), .z (z[1]));
  CDN_mux6 g3(.sel0 (ctl[5]), .data0 (in_0[0]), .sel1 (ctl[4]), .data1
       (in_1[0]), .sel2 (ctl[3]), .data2 (in_2[0]), .sel3 (ctl[2]),
       .data3 (in_3[0]), .sel4 (ctl[1]), .data4 (in_4[0]), .sel5
       (ctl[0]), .data5 (in_5[0]), .z (z[0]));
endmodule

module fx68k_bmux_1464(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     z);
  input [2:0] ctl;
  input [7:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [7:0] z;
  wire [2:0] ctl;
  wire [7:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [7:0] z;
  CDN_bmux7 g1(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .z (z[7]));
  CDN_bmux7 g2(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .z (z[6]));
  CDN_bmux7 g3(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .z (z[5]));
  CDN_bmux7 g4(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .z (z[4]));
  CDN_bmux7 g5(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .z (z[3]));
  CDN_bmux7 g6(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .z (z[2]));
  CDN_bmux7 g7(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .z (z[1]));
  CDN_bmux7 g8(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .z (z[0]));
endmodule

module fx68k_case_box_398(in_0, out_0);
  input [5:0] in_0;
  output [3:0] out_0;
  wire [5:0] in_0;
  wire [3:0] out_0;
  wire n_7, n_8, n_15, n_21, n_23, n_24, n_47;
  not g19 (n_24, in_0[2]);
  nand g1 (n_8, in_0[5], in_0[4], in_0[3], n_24);
  nand g2 (n_7, in_0[1], n_47);
  nor g3 (out_0[3], n_7, n_8);
  nand g5 (n_15, in_0[1], in_0[0]);
  nor g6 (out_0[2], n_15, n_8);
  nand g8 (n_23, n_21, in_0[0]);
  nor g9 (out_0[1], n_23, n_8);
  nor g10 (out_0[0], out_0[3], out_0[2], out_0[1]);
  not g11 (n_47, in_0[0]);
  not g12 (n_21, in_0[1]);
endmodule

module fx68k_mux_1465(ctl, in_0, in_1, in_2, z);
  input [2:0] ctl;
  input [9:0] in_0, in_1, in_2;
  output [9:0] z;
  wire [2:0] ctl;
  wire [9:0] in_0, in_1, in_2;
  wire [9:0] z;
  CDN_mux3 g1(.sel0 (ctl[2]), .data0 (in_0[9]), .sel1 (ctl[1]), .data1
       (in_1[9]), .sel2 (ctl[0]), .data2 (in_2[9]), .z (z[9]));
  CDN_mux3 g11(.sel0 (ctl[2]), .data0 (in_0[8]), .sel1 (ctl[1]), .data1
       (in_1[8]), .sel2 (ctl[0]), .data2 (in_2[8]), .z (z[8]));
  CDN_mux3 g12(.sel0 (ctl[2]), .data0 (in_0[7]), .sel1 (ctl[1]), .data1
       (in_1[7]), .sel2 (ctl[0]), .data2 (in_2[7]), .z (z[7]));
  CDN_mux3 g13(.sel0 (ctl[2]), .data0 (in_0[6]), .sel1 (ctl[1]), .data1
       (in_1[6]), .sel2 (ctl[0]), .data2 (in_2[6]), .z (z[6]));
  CDN_mux3 g14(.sel0 (ctl[2]), .data0 (in_0[5]), .sel1 (ctl[1]), .data1
       (in_1[5]), .sel2 (ctl[0]), .data2 (in_2[5]), .z (z[5]));
  CDN_mux3 g15(.sel0 (ctl[2]), .data0 (in_0[4]), .sel1 (ctl[1]), .data1
       (in_1[4]), .sel2 (ctl[0]), .data2 (in_2[4]), .z (z[4]));
  CDN_mux3 g16(.sel0 (ctl[2]), .data0 (in_0[3]), .sel1 (ctl[1]), .data1
       (in_1[3]), .sel2 (ctl[0]), .data2 (in_2[3]), .z (z[3]));
  CDN_mux3 g17(.sel0 (ctl[2]), .data0 (in_0[2]), .sel1 (ctl[1]), .data1
       (in_1[2]), .sel2 (ctl[0]), .data2 (in_2[2]), .z (z[2]));
  CDN_mux3 g18(.sel0 (ctl[2]), .data0 (in_0[1]), .sel1 (ctl[1]), .data1
       (in_1[1]), .sel2 (ctl[0]), .data2 (in_2[1]), .z (z[1]));
  CDN_mux3 g19(.sel0 (ctl[2]), .data0 (in_0[0]), .sel1 (ctl[1]), .data1
       (in_1[0]), .sel2 (ctl[0]), .data2 (in_2[0]), .z (z[0]));
endmodule

module fx68k_bmux_1502(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [2:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [9:0] z;
  wire [2:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [9:0] z;
  CDN_bmux8 g1(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .sel2
       (ctl[2]), .data4 (in_4[9]), .data5 (in_5[9]), .data6 (in_6[9]),
       .data7 (in_7[9]), .z (z[9]));
  CDN_bmux8 g2(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .sel2
       (ctl[2]), .data4 (in_4[8]), .data5 (in_5[8]), .data6 (in_6[8]),
       .data7 (in_7[8]), .z (z[8]));
  CDN_bmux8 g3(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .data7 (in_7[7]), .z (z[7]));
  CDN_bmux8 g4(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .data7 (in_7[6]), .z (z[6]));
  CDN_bmux8 g5(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .data7 (in_7[5]), .z (z[5]));
  CDN_bmux8 g6(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .data7 (in_7[4]), .z (z[4]));
  CDN_bmux8 g7(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .z (z[3]));
  CDN_bmux8 g8(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .z (z[2]));
  CDN_bmux8 g9(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .z (z[1]));
  CDN_bmux8 g10(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_bmux_1503(ctl, in_0, in_1, z);
  input ctl, in_0, in_1;
  output z;
  wire ctl, in_0, in_1;
  wire z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0), .data1 (in_1), .z (z));
endmodule

module fx68k_bmux_1504(ctl, in_0, in_1, z);
  input ctl;
  input [3:0] in_0, in_1;
  output [3:0] z;
  wire ctl;
  wire [3:0] in_0, in_1;
  wire [3:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_bmux_1505(ctl, in_0, in_1, z);
  input ctl;
  input [5:0] in_0, in_1;
  output [5:0] z;
  wire ctl;
  wire [5:0] in_0, in_1;
  wire [5:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_case_box_404(in_0, out_0);
  input [3:0] in_0;
  output [7:0] out_0;
  wire [3:0] in_0;
  wire [7:0] out_0;
  wire n_5, n_8, n_9, n_11, n_13, n_14, n_15, n_17;
  wire n_21, n_23, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_69, n_70;
  nor g1 (out_0[7], n_5, n_9);
  nand g2 (n_5, n_69, n_70);
  not g3 (n_69, in_0[2]);
  not g4 (n_70, in_0[3]);
  nand g5 (n_9, in_0[1], n_8);
  not g6 (n_8, in_0[0]);
  nor g7 (out_0[6], n_5, n_11);
  nand g8 (n_11, in_0[1], in_0[0]);
  nor g9 (out_0[5], n_13, n_15);
  nand g10 (n_13, in_0[2], n_70);
  nand g11 (n_15, n_14, n_8);
  not g12 (n_14, in_0[1]);
  nor g13 (out_0[4], n_13, n_17);
  nand g14 (n_17, n_14, in_0[0]);
  nor g15 (out_0[3], n_13, n_9);
  nor g16 (out_0[2], n_13, n_11);
  nor g17 (out_0[1], n_15, n_21);
  nand g18 (n_21, n_69, in_0[3]);
  nand g19 (out_0[0], n_28, n_29);
  nand g20 (n_28, n_26, n_27);
  nand g21 (n_26, n_14, n_25);
  and g22 (n_23, in_0[2], n_70);
  and g23 (n_24, n_69, in_0[3]);
  or g24 (n_25, n_23, n_24);
  nand g25 (n_27, in_0[1], n_70);
  nand g26 (n_29, in_0[0], in_0[3]);
endmodule

module fx68k_bmux_1520(ctl, in_0, in_1, z);
  input ctl;
  input [1:0] in_0, in_1;
  output [1:0] z;
  wire ctl;
  wire [1:0] in_0, in_1;
  wire [1:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_mux_1522(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input [2:0] in_0, in_1;
  output [2:0] z;
  wire [1:0] ctl;
  wire [2:0] in_0, in_1;
  wire [2:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[2]), .sel1 (ctl[0]), .data1
       (in_1[2]), .z (z[2]));
  CDN_mux2 g4(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g5(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_mux_1526(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output z;
  wire [7:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0), .sel1 (ctl[6]), .data1
       (in_1), .sel2 (ctl[5]), .data2 (in_2), .sel3 (ctl[4]), .data3
       (in_3), .sel4 (ctl[3]), .data4 (in_4), .sel5 (ctl[2]), .data5
       (in_5), .sel6 (ctl[1]), .data6 (in_6), .sel7 (ctl[0]), .data7
       (in_7), .z (z));
endmodule

module fx68k_mux_1527(ctl, in_0, in_1, in_2, z);
  input [2:0] ctl;
  input in_0, in_1, in_2;
  output z;
  wire [2:0] ctl;
  wire in_0, in_1, in_2;
  wire z;
  CDN_mux3 g1(.sel0 (ctl[2]), .data0 (in_0), .sel1 (ctl[1]), .data1
       (in_1), .sel2 (ctl[0]), .data2 (in_2), .z (z));
endmodule

module fx68k_mux_1529(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, z);
  input [12:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9,
       in_10, in_11, in_12;
  output z;
  wire [12:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9,
       in_10, in_11, in_12;
  wire z;
  CDN_mux13 g1(.sel0 (ctl[12]), .data0 (in_0), .sel1 (ctl[11]), .data1
       (in_1), .sel2 (ctl[10]), .data2 (in_2), .sel3 (ctl[9]), .data3
       (in_3), .sel4 (ctl[8]), .data4 (in_4), .sel5 (ctl[7]), .data5
       (in_5), .sel6 (ctl[6]), .data6 (in_6), .sel7 (ctl[5]), .data7
       (in_7), .sel8 (ctl[4]), .data8 (in_8), .sel9 (ctl[3]), .data9
       (in_9), .sel10 (ctl[2]), .data10 (in_10), .sel11 (ctl[1]),
       .data11 (in_11), .sel12 (ctl[0]), .data12 (in_12), .z (z));
endmodule

module fx68k_mux_1550(ctl, in_0, in_1, in_2, in_3, in_4, z);
  input [4:0] ctl;
  input in_0, in_1, in_2, in_3, in_4;
  output z;
  wire [4:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4;
  wire z;
  CDN_mux5 g1(.sel0 (ctl[4]), .data0 (in_0), .sel1 (ctl[3]), .data1
       (in_1), .sel2 (ctl[2]), .data2 (in_2), .sel3 (ctl[1]), .data3
       (in_3), .sel4 (ctl[0]), .data4 (in_4), .z (z));
endmodule

module fx68k_mux_1577(ctl, in_0, in_1, in_2, in_3, z);
  input [3:0] ctl;
  input in_0, in_1, in_2, in_3;
  output z;
  wire [3:0] ctl;
  wire in_0, in_1, in_2, in_3;
  wire z;
  CDN_mux4 g1(.sel0 (ctl[3]), .data0 (in_0), .sel1 (ctl[2]), .data1
       (in_1), .sel2 (ctl[1]), .data2 (in_2), .sel3 (ctl[0]), .data3
       (in_3), .z (z));
endmodule

module fx68k_mux_1580(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9,
       in_10, in_11;
  output z;
  wire [11:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9,
       in_10, in_11;
  wire z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0), .sel1 (ctl[10]), .data1
       (in_1), .sel2 (ctl[9]), .data2 (in_2), .sel3 (ctl[8]), .data3
       (in_3), .sel4 (ctl[7]), .data4 (in_4), .sel5 (ctl[6]), .data5
       (in_5), .sel6 (ctl[5]), .data6 (in_6), .sel7 (ctl[4]), .data7
       (in_7), .sel8 (ctl[3]), .data8 (in_8), .sel9 (ctl[2]), .data9
       (in_9), .sel10 (ctl[1]), .data10 (in_10), .sel11 (ctl[0]),
       .data11 (in_11), .z (z));
endmodule

module fx68k_bmux_1590(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, z);
  input [3:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9,
       in_10, in_11, in_12, in_13, in_14, in_15;
  output z;
  wire [3:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9,
       in_10, in_11, in_12, in_13, in_14, in_15;
  wire z;
  CDN_bmux16 g1(.sel0 (ctl[0]), .data0 (in_0), .data1 (in_1), .sel1
       (ctl[1]), .data2 (in_2), .data3 (in_3), .sel2 (ctl[2]), .data4
       (in_4), .data5 (in_5), .data6 (in_6), .data7 (in_7), .sel3
       (ctl[3]), .data8 (in_8), .data9 (in_9), .data10 (in_10), .data11
       (in_11), .data12 (in_12), .data13 (in_13), .data14 (in_14),
       .data15 (in_15), .z (z));
endmodule

module fx68k_mux_1611(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, z);
  input [9:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9;
  output z;
  wire [9:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9;
  wire z;
  CDN_mux10 g1(.sel0 (ctl[9]), .data0 (in_0), .sel1 (ctl[8]), .data1
       (in_1), .sel2 (ctl[7]), .data2 (in_2), .sel3 (ctl[6]), .data3
       (in_3), .sel4 (ctl[5]), .data4 (in_4), .sel5 (ctl[4]), .data5
       (in_5), .sel6 (ctl[3]), .data6 (in_6), .sel7 (ctl[2]), .data7
       (in_7), .sel8 (ctl[1]), .data8 (in_8), .sel9 (ctl[0]), .data9
       (in_9), .z (z));
endmodule

module fx68k_bmux_1619(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [2:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output z;
  wire [2:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire z;
  CDN_bmux8 g1(.sel0 (ctl[0]), .data0 (in_0), .data1 (in_1), .sel1
       (ctl[1]), .data2 (in_2), .data3 (in_3), .sel2 (ctl[2]), .data4
       (in_4), .data5 (in_5), .data6 (in_6), .data7 (in_7), .z (z));
endmodule

module fx68k_pla_lined(movEa, col, opcode, lineBmap, palIll, plaA1,
     plaA2, plaA3);
  input [3:0] movEa, col;
  input [15:0] opcode, lineBmap;
  output palIll;
  output [9:0] plaA1, plaA2, plaA3;
  wire [3:0] movEa, col;
  wire [15:0] opcode, lineBmap;
  wire palIll;
  wire [9:0] plaA1, plaA2, plaA3;
  wire [29:0] \cmbsop_arA1[0] ;
  wire [9:0] scA3;
  wire [9:0] \arA23[0] ;
  wire [19:0] \cmbsop_arA1[1] ;
  wire [9:0] \arA23[1] ;
  wire [19:0] \cmbsop_arA1[2] ;
  wire [9:0] \arA23[2] ;
  wire [19:0] \cmbsop_arA1[3] ;
  wire [9:0] \arA23[3] ;
  wire [19:0] \cmbsop_arA1[4] ;
  wire [9:0] \arA23[4] ;
  wire [19:0] \cmbsop_arA1[5] ;
  wire [9:0] \arA23[5] ;
  wire [19:0] \cmbsop_arA1[8] ;
  wire [9:0] \arA23[8] ;
  wire [19:0] \cmbsop_arA1[9] ;
  wire [9:0] \arA23[9] ;
  wire [19:0] \cmbsop_arA1[11] ;
  wire [9:0] \arA23[11] ;
  wire [19:0] \cmbsop_arA1[12] ;
  wire [9:0] \arA23[12] ;
  wire [19:0] \cmbsop_arA1[13] ;
  wire [9:0] \arA23[13] ;
  wire [9:0] \arA23[line] ;
  wire [9:0] \arA1[0] ;
  wire [9:0] \arA1[1] ;
  wire [9:0] \arA1[2] ;
  wire [9:0] \arA1[3] ;
  wire [10:0] cmbsop_a1Misc;
  wire [9:0] a1Misc;
  wire [9:0] \arA1[4] ;
  wire [9:0] \arA1[5] ;
  wire [9:0] \arA1[6] ;
  wire [9:0] \arA1[8] ;
  wire [9:0] \arA1[9] ;
  wire [9:0] \arA1[11] ;
  wire [9:0] \arA1[12] ;
  wire [9:0] \arA1[13] ;
  wire [9:0] \arA1[14] ;
  wire [15:0] arIll;
  wire UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3,
       UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, UNCONNECTED7;
  wire UNCONNECTED8, UNCONNECTED9, UNCONNECTED10, UNCONNECTED11,
       UNCONNECTED12, UNCONNECTED13, UNCONNECTED14, UNCONNECTED15;
  wire UNCONNECTED16, UNCONNECTED17, UNCONNECTED18, UNCONNECTED19,
       UNCONNECTED20, UNCONNECTED21, UNCONNECTED22, UNCONNECTED23;
  wire UNCONNECTED24, UNCONNECTED25, UNCONNECTED26, UNCONNECTED27,
       UNCONNECTED28, UNCONNECTED29, UNCONNECTED30, UNCONNECTED31;
  wire UNCONNECTED32, UNCONNECTED33, UNCONNECTED34, UNCONNECTED35,
       UNCONNECTED36, UNCONNECTED37, UNCONNECTED38, UNCONNECTED39;
  wire UNCONNECTED40, UNCONNECTED41, UNCONNECTED42, UNCONNECTED43,
       UNCONNECTED44, UNCONNECTED45, UNCONNECTED46, UNCONNECTED47;
  wire UNCONNECTED48, UNCONNECTED49, UNCONNECTED50, UNCONNECTED51,
       UNCONNECTED52, UNCONNECTED53, UNCONNECTED54, UNCONNECTED55;
  wire UNCONNECTED56, UNCONNECTED57, UNCONNECTED58, UNCONNECTED59,
       UNCONNECTED60, UNCONNECTED61, UNCONNECTED62, UNCONNECTED63;
  wire UNCONNECTED64, UNCONNECTED65, UNCONNECTED66, UNCONNECTED67,
       UNCONNECTED68, UNCONNECTED69, UNCONNECTED70, UNCONNECTED71;
  wire UNCONNECTED72, UNCONNECTED73, UNCONNECTED74, UNCONNECTED75,
       UNCONNECTED76, UNCONNECTED77, UNCONNECTED78, UNCONNECTED79;
  wire UNCONNECTED80, UNCONNECTED81, UNCONNECTED82, UNCONNECTED83,
       UNCONNECTED84, UNCONNECTED85, UNCONNECTED86, UNCONNECTED87;
  wire UNCONNECTED88, UNCONNECTED89, UNCONNECTED90, UNCONNECTED91,
       UNCONNECTED92, UNCONNECTED93, UNCONNECTED94, UNCONNECTED95;
  wire UNCONNECTED96, UNCONNECTED97, UNCONNECTED98, UNCONNECTED99,
       UNCONNECTED100, UNCONNECTED101, UNCONNECTED102, UNCONNECTED103;
  wire UNCONNECTED104, UNCONNECTED105, UNCONNECTED106, UNCONNECTED107,
       UNCONNECTED108, UNCONNECTED109, UNCONNECTED110, UNCONNECTED111;
  wire UNCONNECTED112, UNCONNECTED113, UNCONNECTED114, UNCONNECTED115,
       UNCONNECTED116, UNCONNECTED117, UNCONNECTED118, UNCONNECTED119;
  wire UNCONNECTED120, UNCONNECTED121, UNCONNECTED122, UNCONNECTED123,
       UNCONNECTED124, UNCONNECTED125, UNCONNECTED126, UNCONNECTED127;
  wire UNCONNECTED128, UNCONNECTED129, UNCONNECTED130, UNCONNECTED131,
       UNCONNECTED132, UNCONNECTED133, UNCONNECTED134, UNCONNECTED135;
  wire UNCONNECTED136, UNCONNECTED137, UNCONNECTED138, UNCONNECTED139,
       UNCONNECTED140, UNCONNECTED141, UNCONNECTED142, UNCONNECTED143;
  wire UNCONNECTED144, UNCONNECTED145, UNCONNECTED146, UNCONNECTED147,
       UNCONNECTED148, UNCONNECTED149, UNCONNECTED150, UNCONNECTED151;
  wire UNCONNECTED152, UNCONNECTED153, UNCONNECTED154, UNCONNECTED155,
       UNCONNECTED156, UNCONNECTED157, UNCONNECTED158, UNCONNECTED159;
  wire UNCONNECTED160, UNCONNECTED161, UNCONNECTED162, UNCONNECTED163,
       UNCONNECTED164, UNCONNECTED165, UNCONNECTED166, UNCONNECTED167;
  wire UNCONNECTED168, UNCONNECTED169, UNCONNECTED170, UNCONNECTED171,
       UNCONNECTED172, UNCONNECTED173, UNCONNECTED174, UNCONNECTED175;
  wire UNCONNECTED176, UNCONNECTED177, UNCONNECTED178, UNCONNECTED179,
       UNCONNECTED180, UNCONNECTED181, UNCONNECTED182, UNCONNECTED183;
  wire UNCONNECTED184, UNCONNECTED185, UNCONNECTED186, UNCONNECTED187,
       UNCONNECTED188, UNCONNECTED189, UNCONNECTED190, UNCONNECTED191;
  wire UNCONNECTED192, UNCONNECTED193, UNCONNECTED194, UNCONNECTED195,
       UNCONNECTED196, UNCONNECTED197, UNCONNECTED198, UNCONNECTED199;
  wire UNCONNECTED200, UNCONNECTED201, UNCONNECTED202, UNCONNECTED203,
       UNCONNECTED204, UNCONNECTED205, UNCONNECTED206, UNCONNECTED207;
  wire UNCONNECTED208, UNCONNECTED209, UNCONNECTED210, UNCONNECTED211,
       UNCONNECTED212, UNCONNECTED213, UNCONNECTED214, UNCONNECTED215;
  wire UNCONNECTED216, UNCONNECTED217, UNCONNECTED218, UNCONNECTED219,
       UNCONNECTED220, UNCONNECTED221, UNCONNECTED222, UNCONNECTED223;
  wire UNCONNECTED224, UNCONNECTED225, UNCONNECTED226, UNCONNECTED227,
       UNCONNECTED228, UNCONNECTED229, UNCONNECTED230, UNCONNECTED231;
  wire UNCONNECTED232, UNCONNECTED233, UNCONNECTED234, UNCONNECTED235,
       UNCONNECTED236, UNCONNECTED237, UNCONNECTED238, UNCONNECTED239;
  wire UNCONNECTED240, UNCONNECTED241, UNCONNECTED242, UNCONNECTED243,
       UNCONNECTED244, UNCONNECTED245, UNCONNECTED246, UNCONNECTED247;
  wire UNCONNECTED248, UNCONNECTED249, UNCONNECTED250, UNCONNECTED251,
       UNCONNECTED252, UNCONNECTED253, UNCONNECTED254, UNCONNECTED255;
  wire UNCONNECTED256, UNCONNECTED257, UNCONNECTED258, UNCONNECTED259,
       UNCONNECTED260, UNCONNECTED261, UNCONNECTED262, UNCONNECTED263;
  wire UNCONNECTED264, UNCONNECTED265, UNCONNECTED266, UNCONNECTED267,
       UNCONNECTED268, UNCONNECTED269, UNCONNECTED270, UNCONNECTED271;
  wire UNCONNECTED272, UNCONNECTED273, UNCONNECTED274, UNCONNECTED275,
       UNCONNECTED276, UNCONNECTED277, UNCONNECTED278, UNCONNECTED279;
  wire UNCONNECTED280, UNCONNECTED281, UNCONNECTED282, UNCONNECTED283,
       UNCONNECTED284, UNCONNECTED285, UNCONNECTED286, UNCONNECTED287;
  wire UNCONNECTED288, UNCONNECTED289, UNCONNECTED290, UNCONNECTED291,
       UNCONNECTED292, UNCONNECTED293, UNCONNECTED294, UNCONNECTED295;
  wire UNCONNECTED296, UNCONNECTED297, UNCONNECTED298, UNCONNECTED299,
       UNCONNECTED300, UNCONNECTED301, UNCONNECTED302, UNCONNECTED303;
  wire UNCONNECTED304, UNCONNECTED305, UNCONNECTED306, UNCONNECTED307,
       UNCONNECTED308, UNCONNECTED309, UNCONNECTED310, UNCONNECTED311;
  wire UNCONNECTED312, UNCONNECTED313, UNCONNECTED314, UNCONNECTED315,
       UNCONNECTED316, UNCONNECTED317, UNCONNECTED318, UNCONNECTED319;
  wire UNCONNECTED320, UNCONNECTED321, UNCONNECTED322, UNCONNECTED323,
       UNCONNECTED324, UNCONNECTED325, UNCONNECTED326, UNCONNECTED327;
  wire UNCONNECTED328, UNCONNECTED329, UNCONNECTED330, UNCONNECTED331,
       UNCONNECTED332, UNCONNECTED333, UNCONNECTED334, UNCONNECTED335;
  wire UNCONNECTED336, UNCONNECTED337, UNCONNECTED338, UNCONNECTED339,
       UNCONNECTED340, UNCONNECTED341, UNCONNECTED342, UNCONNECTED343;
  wire UNCONNECTED344, UNCONNECTED345, UNCONNECTED346, UNCONNECTED347,
       UNCONNECTED348, UNCONNECTED349, UNCONNECTED350, UNCONNECTED351;
  wire UNCONNECTED352, UNCONNECTED353, UNCONNECTED354, UNCONNECTED355,
       UNCONNECTED356, UNCONNECTED357, UNCONNECTED358, UNCONNECTED359;
  wire UNCONNECTED360, UNCONNECTED361, UNCONNECTED362, UNCONNECTED363,
       UNCONNECTED364, UNCONNECTED365, UNCONNECTED366, UNCONNECTED367;
  wire UNCONNECTED368, UNCONNECTED369, UNCONNECTED370, UNCONNECTED371,
       UNCONNECTED372, UNCONNECTED373, UNCONNECTED374, UNCONNECTED375;
  wire UNCONNECTED376, UNCONNECTED377, UNCONNECTED378, UNCONNECTED379,
       UNCONNECTED380, UNCONNECTED381, UNCONNECTED382, UNCONNECTED383;
  wire UNCONNECTED384, UNCONNECTED385, UNCONNECTED386, UNCONNECTED387,
       UNCONNECTED388, UNCONNECTED389, UNCONNECTED390, UNCONNECTED391;
  wire UNCONNECTED392, UNCONNECTED393, UNCONNECTED394, UNCONNECTED395,
       UNCONNECTED396, UNCONNECTED397, UNCONNECTED398, UNCONNECTED399;
  wire UNCONNECTED400, UNCONNECTED401, UNCONNECTED402, UNCONNECTED403,
       UNCONNECTED404, UNCONNECTED405, UNCONNECTED406, UNCONNECTED407;
  wire UNCONNECTED408, UNCONNECTED409, UNCONNECTED410, UNCONNECTED411,
       UNCONNECTED412, UNCONNECTED413, UNCONNECTED414, UNCONNECTED415;
  wire UNCONNECTED416, UNCONNECTED417, UNCONNECTED418, UNCONNECTED419,
       UNCONNECTED420, UNCONNECTED421, UNCONNECTED422, UNCONNECTED423;
  wire UNCONNECTED424, _X_, illMisc, n_7, n_8, n_10, n_14, n_15;
  wire n_17, n_19, n_22, n_23, n_24, n_26, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_40, n_41, n_43, n_44;
  wire n_46, n_47, n_48, n_64, n_67, n_73, n_79, n_81;
  wire n_82, n_83, n_87, n_88, n_101, n_114, n_124, n_125;
  wire n_152, n_153, n_154, n_167, n_23477, n_23482, n_23483, n_23484;
  wire n_23485, n_23486, n_23487, n_23488, n_23489, n_23490, n_23491,
       n_23492;
  wire n_23493, n_23494, n_23495, n_23496, n_23497, n_23498, n_23499,
       n_23500;
  wire n_23501, n_23502, n_23503, n_23504, n_23505, n_23506, n_23507,
       n_23508;
  wire n_23509, n_23510, n_23511, n_23512, n_23513, n_23514, n_23515,
       n_23516;
  wire n_23517, n_23518, n_23519, n_23520, n_23521, n_23522, n_23523,
       n_23524;
  wire n_23525, n_23526, n_23527, n_23528, n_23529, n_23530, n_23531,
       n_23532;
  wire n_23533, n_23534, n_23535, n_23536, n_23537, n_23538, n_23539,
       n_23540;
  wire n_23541, n_23542, n_23543, n_23544, n_23545, n_23546, n_23547,
       n_23548;
  wire n_23549, n_23550, n_23551, n_23552, n_23553, n_23554, n_23555,
       n_23556;
  wire n_23557, n_23558, n_23559, n_23560, n_23561, n_23562, n_23563,
       n_23564;
  wire n_23565, n_23566, n_23567, n_23568, n_23569, n_23570, n_23571,
       n_23572;
  wire n_23573, n_23574, n_23575, n_23576, n_23577, n_23578, n_23579,
       n_23580;
  wire n_23581, n_23582, n_23583, n_23584, n_23585, n_23586, n_23587,
       n_23588;
  wire n_23589, n_23590, n_23591, n_23592, n_23593, n_23594, n_23595,
       n_23596;
  wire n_23597, n_23598, n_23599, n_23600, n_23601, n_23602, n_23603,
       n_23604;
  wire n_23605, n_23606, n_23607, n_23608, n_23609, n_23610, n_23611,
       n_23612;
  wire n_23613, n_23614, n_23615, n_23616, n_23617, n_23618, n_23619,
       n_23620;
  wire n_23621, n_23622, n_23623, n_23624, n_23625, n_23626, n_23627,
       n_23628;
  wire n_23629, n_23630, n_23631, n_23632, n_23633, n_23634, n_23635,
       n_23636;
  wire n_23637, n_23638, n_23639, n_23640, n_23641, n_23642, n_23643,
       n_23644;
  wire n_23645, n_23646, n_23647, n_23648, n_23649, n_23650, n_23651,
       n_23652;
  wire n_23653, n_23654, n_23655, n_23656, n_23657, n_23658, n_23665,
       n_23666;
  wire n_23667, n_23668, n_23669, n_23670, n_23671, n_23682, n_23683,
       n_23684;
  wire n_23685, n_23686, n_23687, n_23688, n_23689, n_23690, n_23697,
       n_23698;
  wire n_23699, n_23700, n_23701, n_23702, n_23703, n_23704, n_23705,
       n_23706;
  wire n_23707, n_23708, n_23709, n_23710, n_23711, n_23712, n_23713,
       n_23714;
  wire n_23715, n_23716, n_23717, n_23718, n_23719, n_23720, n_23721,
       n_23722;
  wire n_23723, n_23724, n_23725, n_23726, n_23727, n_23728, n_23729,
       n_23730;
  wire n_23731, n_23732, n_23733, n_23734, n_23735, n_23736, n_23737,
       n_23738;
  wire n_23739, n_23740, n_23741, n_23742, n_23743, n_23744, n_23745,
       n_23746;
  wire n_23747, n_23748, n_23749, n_23750, n_23751, n_23752, n_23753,
       n_23754;
  wire n_23755, n_23756, n_23757, n_23758, n_23759, n_23760, n_23761,
       n_23762;
  wire n_23763, n_23764, n_23765, n_23766, n_23767, n_23768, n_23769,
       n_23770;
  wire n_23771, n_23772, n_23773, n_23774, n_23775, n_23776, n_23777,
       n_23778;
  wire n_23779, n_23780, n_23781, n_23782, n_23783, n_23784, n_23785,
       n_23786;
  wire n_23787, n_23788, n_23789, n_23790, n_23791, n_23792, n_23793,
       n_23794;
  wire n_23795, n_23796, n_23797, n_23798, n_23799, n_23800, n_23801,
       n_23802;
  wire n_23803, n_23804, n_23805, n_23806, n_23807, n_23808, n_23809,
       n_23810;
  wire n_23811, n_23812, n_23813, n_23814, n_23815, n_23816, n_23817,
       n_23818;
  wire n_23819, n_23820, n_23821, n_23822, n_23823, n_23824, n_23825,
       n_23826;
  wire n_23827, n_23828, n_23829, n_23830, n_23831, n_23832, n_23833,
       n_23834;
  wire n_23835, n_23836, n_23837, n_23838, n_23839, n_23840, n_23841,
       n_23842;
  wire n_23843, n_23844, n_23845, n_23846, n_23847, n_23848, n_23849,
       n_23850;
  wire n_23851, n_23852, n_23853, n_23854, n_23855, n_23856, n_23857,
       n_23858;
  wire n_23859, n_23860, n_23861, n_23862, n_23863, n_23864, n_23865,
       n_23866;
  wire n_23867, n_23868, n_23869, n_23870, n_23871, n_23872, n_23873,
       n_23874;
  wire n_23875, n_23876, n_23877, n_23878, n_23879, n_23880, n_23881,
       n_23882;
  wire n_23883, n_23884, n_23885, n_23886, n_23887, n_23888, n_23889,
       n_23890;
  wire n_23891, n_23892, n_23893, n_23894, n_23895, n_23896, n_23897,
       n_23898;
  wire n_23899, n_23900, n_23901, n_23902, n_23903, n_23904, n_23905,
       n_23906;
  wire n_23907, n_23908, n_23909, n_23910, n_23911, n_23912, n_23913,
       n_23914;
  wire n_23915, n_23916, n_23917, n_23918, n_23919, n_23920, n_23921,
       n_23922;
  wire n_23923, n_23924, n_23925, n_23926, n_23927, n_23928, n_23929,
       n_23930;
  wire n_23931, n_23932, n_23933, n_23934, n_23935, n_23936, n_23937,
       n_23938;
  wire n_23939, n_23940, n_23941, n_23942, n_23943, n_23944, n_23945,
       n_23946;
  wire n_23947, n_23948, n_23949, n_23950, n_23951, n_23952, n_23953,
       n_23954;
  wire n_23955, n_23956, n_23957, n_23958, n_23959, n_23960, n_23961,
       n_23962;
  wire n_23963, n_23964, n_23965, n_23966, n_23967, n_23968, n_23969,
       n_23970;
  wire n_23971, n_23972, n_23973, n_23974, n_23975, n_23976, n_23977,
       n_23978;
  wire n_23979, n_23980, n_23981, n_23982, n_23983, n_23984, n_23985,
       n_23986;
  wire n_23987, n_23988, n_23989, n_23990, n_23991, n_23992, n_23993,
       n_23994;
  wire n_23995, n_23996, n_23997, n_23998, n_23999, n_24000, n_24001,
       n_24002;
  wire n_24003, n_24004, n_24005, n_24006, n_24007, n_24008, n_24009,
       n_24010;
  wire n_24011, n_24012, n_24013, n_24014, n_24015, n_24016, n_24017,
       n_24018;
  wire n_24019, n_24020, n_24021, n_24022, n_24023, n_24024, n_24025,
       n_24026;
  wire n_24027, n_24028, n_24029, n_24030, n_24031, n_24032, n_24033,
       n_24034;
  wire n_24035, n_24036, n_24037, n_24038, n_24039, n_24040, n_24041,
       n_24042;
  wire n_24043, n_24044, n_24045, n_24046, n_24047, n_24048, n_24049,
       n_24050;
  wire n_24051, n_24052, n_24053, n_24058, n_24059, n_24060, n_24061,
       n_24062;
  wire n_24063, n_24064, n_24065, n_24066, n_24067, n_24068, n_24069,
       n_24070;
  wire n_24071, n_24072, n_24073, n_24074, n_24075, n_24076, n_24077,
       n_24078;
  wire n_24079, n_24080, n_24081, n_24082, n_24083, n_24084, n_24085,
       n_24086;
  wire n_24087, n_24088, n_24089, n_24090, n_24091, n_24092, n_24093,
       n_24094;
  wire n_24095, n_24096, n_24097, n_24098, n_24099, n_24100, n_24101,
       n_24102;
  wire n_24103, n_24104, n_24105, n_24106, n_24107, n_24108, n_24109,
       n_24110;
  wire n_24111, n_24112, n_24113, n_24114, n_24115, n_24116, n_24117,
       n_24118;
  wire n_24119, n_24120, n_24121, n_24122, n_24123, n_24124, n_24125,
       n_24126;
  wire n_24127, n_24128, n_24129, n_24130, n_24131, n_24132, n_24133,
       n_24134;
  wire n_24135, n_24136, n_24137, n_24138, n_24139, n_24140, n_24141,
       n_24142;
  wire n_24143, n_24144, n_24145, n_24146, n_24147, n_24148, n_24149,
       n_24150;
  wire n_24151, n_24152, n_24153, n_24154, n_24155, n_24156, n_24157,
       n_24158;
  wire n_24159, n_24160, n_24161, n_24162, n_24163, n_24164, n_24165,
       n_24166;
  wire n_24167, n_24168, n_24169, n_24170, n_24171, n_24172, n_24173,
       n_24174;
  wire n_24175, n_24176, n_24177, n_24178, n_24179, n_24180, n_24181,
       n_24182;
  wire n_24183, n_24184, n_24185, n_24186, n_24187, n_24188, n_24189,
       n_24190;
  wire n_24191, n_24192, n_24193, n_24194, n_24195, n_24196, n_24197,
       n_24198;
  wire n_24199, n_24200, n_24201, n_24202, n_24203, n_24204, n_24205,
       n_24206;
  wire n_24207, n_24208, n_24209, n_24210, n_24211, n_24212, n_24213,
       n_24214;
  wire n_24215, n_24216, n_24217, n_24218, n_24219, n_24220, n_24221,
       n_24222;
  wire n_24223, n_24224, n_24225, n_24226, n_24227, n_24228, n_24229,
       n_24230;
  wire n_24231, n_24232, n_24233, n_24234, n_24235, n_24236, n_24237,
       n_24238;
  wire n_24239, n_24240, n_24241, n_24242, n_24243, n_24244, n_24245,
       n_24246;
  wire n_24247, n_24248, n_24249, n_24250, n_24251, n_24252, n_24253,
       n_24254;
  wire n_24255, n_24256, n_24257, n_24258, n_24259, n_24260, n_24261,
       n_24262;
  wire n_24263, n_24264, n_24265, n_24266, n_24267, n_24268, n_24269,
       n_24270;
  wire n_24271, n_24272, n_24273, n_24274, n_24275, n_24276, n_24277,
       n_24278;
  wire n_24279, n_24280, n_24281, n_24282, n_24283, n_24284, n_24285,
       n_24286;
  wire n_24287, n_24288, n_24289, n_24290, n_24291, n_24292, n_24293,
       n_24294;
  wire n_24295, n_24296, n_24297, n_24298, n_24299, n_24300, n_24301,
       n_24302;
  wire n_24303, n_24304, n_24305, n_24306, n_24307, n_24308, n_24309,
       n_24310;
  wire n_24311, n_24312, n_24313, n_24314, n_24315, n_24316, n_24317,
       n_24318;
  wire n_24319, n_24320, n_24321, n_24322, n_24323, n_24324, n_24325,
       n_24326;
  wire n_24327, n_24328, n_24329, n_24330, n_24331, n_24332, n_24333,
       n_24334;
  wire n_24335, n_24336, n_24337, n_24338, n_24339, n_24340, n_24341,
       n_24342;
  wire n_24343, n_24344, n_24345, n_24346, n_24347, n_24348, n_24349,
       n_24350;
  wire n_24351, n_24352, n_24353, n_24354, n_24355, n_24356, n_24357,
       n_24358;
  wire n_24359, n_24360, n_24361, n_24362, n_24363, n_24364, n_24365,
       n_24366;
  wire n_24367, n_24368, n_24369, n_24370, n_24371, n_24372, n_24373,
       n_24374;
  wire n_24375, n_24376, n_24377, n_24378, n_24379, n_24380, n_24381,
       n_24382;
  wire n_24383, n_24384, n_24385, n_24386, n_24387, n_24388, n_24389,
       n_24390;
  wire n_24391, n_24392, n_24393, n_24394, n_24395, n_24396, n_24397,
       n_24398;
  wire n_24399, n_24400, n_24401, n_24402, n_24403, n_24404, n_24405,
       n_24406;
  wire n_24407, n_24408, n_24409, n_24410, n_24411, n_24412, n_24413,
       n_24414;
  wire n_24415, n_24416, n_24417, n_24418, n_24419, n_24420, n_24421,
       n_24422;
  wire n_24423, n_24424, n_24425, n_24426, n_24427, n_24428, n_24429,
       n_24430;
  wire n_24431, n_24432, n_24433, n_24434, n_24435, n_24436, n_24437,
       n_24438;
  wire n_24439, n_24440, n_24441, n_24442, n_24443, n_24444, n_24445,
       n_24446;
  wire n_24447, n_24448, n_24449, n_24450, n_24451, n_24452, n_24453,
       n_24454;
  wire n_24455, n_24456, n_24457, n_24458, n_24459, n_24460, n_24461,
       n_24462;
  wire n_24463, n_24464, n_24465, n_24466, n_24467, n_24468, n_24469,
       n_24470;
  wire n_24471, n_24472, n_24473, n_24474, n_24475, n_24476, n_24477,
       n_24478;
  wire n_24479, n_24480, n_24481, n_24482, n_24483, n_24484, n_24485,
       n_24486;
  wire n_24487, n_24488, n_24489, n_24490, n_24491, n_24492, n_24493,
       n_24494;
  wire n_24495, n_24496, n_24497, n_24498, n_24499, n_24500, n_24501,
       n_24502;
  wire n_24503, n_24504, n_24505, n_24506, n_24507, n_24508, n_24509,
       n_24510;
  wire n_24511, n_24512, n_24513, n_24514, n_24515, n_24516, n_24517,
       n_24518;
  wire n_24519, n_24520, n_24521, n_24522, n_24523, n_24524, n_24525,
       n_24526;
  wire n_24527, n_24528, n_24529, n_24536, n_24537, n_24538, n_24539,
       n_24540;
  wire n_24541, n_24542, n_24543, n_24544, n_24545, n_24546, n_24547,
       n_24548;
  wire n_24549, n_24550, n_24551, n_24552, n_24553, n_24554, n_24555,
       n_24556;
  wire n_24557, n_24558, n_24559, n_24560, n_24561, n_24562, n_24563,
       n_24564;
  wire n_24565, n_24566, n_24567, n_24568, n_24569, n_24570, n_24571,
       n_24572;
  wire n_24573, n_24574, n_24575, n_24576, n_24577, n_24578, n_24579,
       n_24580;
  wire n_24581, n_24582, n_24583, n_24584, n_24585, n_24586, n_24587,
       n_24588;
  wire n_24589, n_24590, n_24591, n_24592, n_24593, n_24594, n_24595,
       n_24596;
  wire n_24597, n_24598, n_24599, n_24600, n_24601, n_24602, n_24603,
       n_24604;
  wire n_24605, n_24606, n_24607, n_24608, n_24609, n_24610, n_24611,
       n_24612;
  wire n_24613, n_24614, n_24615, n_24616, n_24617, n_24618, n_24619,
       n_24620;
  wire n_24621, n_24622, n_24627, n_24628, n_24629, n_24630, n_24631,
       n_24632;
  wire n_24633, n_24634, n_24635, n_24636, n_24637, n_24638, n_24639,
       n_24640;
  wire n_24641, n_24642, n_24643, n_24644, n_24645, n_24646, n_24647,
       n_24648;
  wire n_24649, n_24650, n_24651, n_24652, n_24653, n_24654, n_24655,
       n_24656;
  wire n_24657, n_24658, n_24659, n_24660, n_24661, n_24662, n_24663,
       n_24664;
  wire n_24665, n_24666, n_24667, n_24668, n_24669, n_24670, n_24671,
       n_24672;
  wire n_24673, n_24674, n_24675, n_24676, n_24677, n_24678, n_24679,
       n_24680;
  wire n_24681, n_24682, n_24683, n_24684, n_24685, n_24686, n_24687,
       n_24688;
  wire n_24689, n_24690, n_24691, n_24692, n_24693, n_24694, n_24695,
       n_24696;
  wire n_24697, n_24698, n_24699, n_24700, n_24701, n_24702, n_24703,
       n_24704;
  wire n_24713, n_24714, n_24715, n_24716, n_24717, n_24718, n_24719,
       n_24720;
  wire n_24721, n_24722, n_24723, n_24724, n_24725, n_24726, n_24727,
       n_24728;
  wire n_24729, n_24730, n_24731, n_24732, n_24733, n_24734, n_24735,
       n_24736;
  wire n_24737, n_24738, n_24739, n_24740, n_24741, n_24742, n_24743,
       n_24744;
  wire n_24745, n_24746, n_24747, n_24748, n_24749, n_24750, n_24751,
       n_24752;
  wire n_24753, n_24754, n_24755, n_24756, n_24757, n_24758, n_24759,
       n_24760;
  wire n_24761, n_24762, n_24763, n_24764, n_24765, n_24766, n_24767,
       n_24768;
  wire n_24769, n_24770, n_24771, n_24772, n_24773, n_24774, n_24775,
       n_24776;
  wire n_24777, n_24778, n_24779, n_24780, n_24781, n_24782, n_24783,
       n_24784;
  wire n_24785, n_24786, n_24787, n_24788, n_24789, n_24790, n_24791,
       n_24792;
  wire n_24793, n_24794, n_24795, n_24796, n_24797, n_24798, n_24799,
       n_24800;
  wire n_24801, n_24802, n_24803, n_24804, n_24813, n_24814, n_24815,
       n_24816;
  wire n_24817, n_24818, n_24819, n_24820, n_24821, n_24822, n_24823,
       n_24824;
  wire n_24825, n_24826, n_24827, n_24828, n_24829, n_24830, n_24831,
       n_24832;
  wire n_24833, n_24834, n_24835, n_24836, n_24837, n_24838, n_24839,
       n_24840;
  wire n_24841, n_24842, n_24843, n_24844, n_24845, n_24846, n_24847,
       n_24848;
  wire n_24849, n_24850, n_24851, n_24852, n_24853, n_24854, n_24855,
       n_24856;
  wire n_24857, n_24858, n_24859, n_24860, n_24861, n_24862, n_24863,
       n_24864;
  wire n_24865, n_24866, n_24867, n_24868, n_24869, n_24870, n_24871,
       n_24872;
  wire n_24873, n_24874, n_24875, n_24876, n_24877, n_24878, n_24879,
       n_24880;
  wire n_24881, n_24882, n_24883, n_24884, n_24885, n_24886, n_24887,
       n_24888;
  wire n_24889, n_24890, n_24891, n_24892, n_24893, n_24894, n_24895,
       n_24896;
  wire n_24897, n_24898, n_24899, n_24900, n_24901, n_24902, n_24903,
       n_24904;
  wire n_24905, n_24906, n_24907, n_24908, n_24917, n_24918, n_24919,
       n_24920;
  wire n_24921, n_24922, n_24923, n_24924, n_24925, n_24926, n_24927,
       n_24928;
  wire n_24929, n_24930, n_24931, n_24932, n_24933, n_24934, n_24935,
       n_24936;
  wire n_24937, n_24938, n_24939, n_24940, n_24941, n_24942, n_24943,
       n_24944;
  wire n_24945, n_24946, n_24947, n_24948, n_24949, n_24950, n_24951,
       n_24952;
  wire n_24953, n_24954, n_24955, n_24956, n_24957, n_24958, n_24959,
       n_24960;
  wire n_24961, n_24962, n_24963, n_24964, n_24965, n_24966, n_24967,
       n_24968;
  wire n_24969, n_24970, n_24971, n_24972, n_24973, n_24974, n_24975,
       n_24976;
  wire n_24977, n_24978, n_24979, n_24980, n_24981, n_24982, n_24983,
       n_24984;
  wire n_24985, n_24986, n_24987, n_24988, n_24989, n_24990, n_24991,
       n_24992;
  wire n_24993, n_24994, n_24995, n_24996, n_24997, n_24998, n_24999,
       n_25000;
  wire n_25001, n_25002, n_25003, n_25012, n_25013, n_25014, n_25015,
       n_25016;
  wire n_25017, n_25018, n_25019, n_25020, n_25021, n_25022, n_25023,
       n_25024;
  wire n_25025, n_25026, n_25027, n_25028, n_25029, n_25030, n_25031,
       n_25032;
  wire n_25033, n_25034, n_25035, n_25036, n_25037, n_25038, n_25039,
       n_25040;
  wire n_25041, n_25042, n_25043, n_25044, n_25045, n_25046, n_25047,
       n_25048;
  wire n_25049, n_25050, n_25051, n_25052, n_25053, n_25054, n_25055,
       n_25056;
  wire n_25057, n_25058, n_25059, n_25060, n_25061, n_25062, n_25063,
       n_25064;
  wire n_25065, n_25066, n_25067, n_25068, n_25069, n_25070, n_25071,
       n_25072;
  wire n_25073, n_25074, n_25075, n_25076, n_25077, n_25078, n_25079,
       n_25080;
  wire n_25081, n_25082, n_25083, n_25084, n_25085, n_25086, n_25087,
       n_25088;
  wire n_25089, n_25090, n_25091, n_25092, n_25093, n_25094, n_25095,
       n_25096;
  wire n_25097, n_25098, n_25099, n_25100, n_25101, n_25102, n_25103,
       n_25112;
  wire n_25113, n_25114, n_25115, n_25116, n_25117, n_25118, n_25119,
       n_25120;
  wire n_25121, n_25122, n_25123, n_25124, n_25125, n_25126, n_25127,
       n_25128;
  wire n_25129, n_25130, n_25131, n_25132, n_25133, n_25134, n_25135,
       n_25136;
  wire n_25137, n_25138, n_25139, n_25140, n_25141, n_25142, n_25143,
       n_25144;
  wire n_25145, n_25146, n_25147, n_25148, n_25149, n_25150, n_25151,
       n_25152;
  wire n_25153, n_25154, n_25155, n_25156, n_25157, n_25158, n_25159,
       n_25160;
  wire n_25161, n_25162, n_25163, n_25164, n_25165, n_25166, n_25167,
       n_25168;
  wire n_25169, n_25170, n_25171, n_25172, n_25173, n_25174, n_25175,
       n_25176;
  wire n_25177, n_25178, n_25179, n_25180, n_25181, n_25182, n_25183,
       n_25184;
  wire n_25185, n_25186, n_25187, n_25188, n_25189, n_25190, n_25191,
       n_25192;
  wire n_25193, n_25194, n_25195, n_25196, n_25197, n_25198, n_25199,
       n_25200;
  wire n_25201, n_25202, n_25203, n_25204, n_25205, n_25206, n_25207,
       n_25208;
  wire n_25209, n_25210, n_25211, n_25212, n_25213, n_25214, n_25215,
       n_25216;
  wire n_25217, n_25218, n_25219, n_25220, n_25221, n_25222, n_25223,
       n_25224;
  wire n_25225, n_25226, n_25227, n_25228, n_25229, n_25230, n_25231,
       n_25232;
  wire n_25233, n_25234, n_25235, n_25236, n_25237, n_25238, n_25239,
       n_25240;
  wire n_25241, n_25242, n_25243, n_25244, n_25245, n_25246, n_25247,
       n_25248;
  wire n_25249, n_25250, n_25251, n_25252, n_25253, n_25254, n_25255,
       n_25256;
  wire n_25257, n_25258, n_25259, n_25260, n_25261, n_25262, n_25263,
       n_25264;
  wire n_25265, n_25266, n_25267, n_25268, n_25269, n_25270, n_25271,
       n_25272;
  wire n_25273, n_25274, n_25275, n_25276, n_25277, n_25278, n_25279,
       n_25280;
  wire n_25281, n_25282, n_25283, n_25284, n_25285, n_25286, n_25287,
       n_25288;
  wire n_25289, n_25290, n_25291, n_25292, n_25293, n_25294, n_25295,
       n_25296;
  wire n_25297, n_25298, n_25299, n_25300, n_25301, n_25302, n_25303,
       n_25304;
  wire n_25305, n_25306, n_25307, n_25308, n_25309, n_25310, n_25311,
       n_25312;
  wire n_25313, n_25314, n_25315, n_25316, n_25317, n_25318, n_25319,
       n_25320;
  wire n_25321, n_25322, n_25323, n_25324, n_25325, n_25326, n_25327,
       n_25328;
  wire n_25329, n_25330, n_25331, n_25332, n_25333, n_25334, n_25335,
       n_25336;
  wire n_25337, n_25338, n_25339, n_25340, n_25341, n_25342, n_25343,
       n_25344;
  wire n_25345, n_25346, n_25347, n_25348, n_25349, n_25350, n_25351,
       n_25352;
  wire n_25353, n_25354, n_25355, n_25356, n_25357, n_25358, n_25359,
       n_25360;
  wire n_25361, n_25362, n_25363, n_25364, n_25365, n_25366, n_25367,
       n_25368;
  wire n_25369, n_25370, n_25371, n_25372, n_25373, n_25374, n_25375,
       n_25376;
  wire n_25377, n_25378, n_25379, n_25380, n_25381, n_25382, n_25383,
       n_25384;
  wire n_25385, n_25386, n_25387, n_25388, n_25389, n_25390, n_25391,
       n_25392;
  wire n_25393, n_25394, n_25395, n_25396, n_25397, n_25398, n_25399,
       n_25400;
  wire n_25401, n_25402, n_25403, n_25404, n_25405, n_25406, n_25407,
       n_25408;
  wire n_25409, n_25410, n_25411, n_25412, n_25413, n_25414, n_25415,
       n_25416;
  wire n_25417, n_25418, n_25419, n_25420, n_25421, n_25422, n_25423,
       n_25424;
  wire n_25425, n_25426, n_25427, n_25428, n_25429, n_25430, n_25431,
       n_25432;
  wire n_25433, n_25434, n_25435, n_25436, n_25437, n_25438, n_25439,
       n_25440;
  wire n_25441, n_25442, n_25443, n_25444, n_25445, n_25446, n_25447,
       n_25448;
  wire n_25449, n_25450, n_25451, n_25452, n_25453, n_25454, n_25455,
       n_25456;
  wire n_25457, n_25458, n_25459, n_25460, n_25461, n_25462, n_25463,
       n_25464;
  wire n_25465, n_25466, n_25467, n_25468, n_25469, n_25470, n_25471,
       n_25472;
  wire n_25473, n_25474, n_25475, n_25476, n_25477, n_25478, n_25479,
       n_25480;
  wire n_25481, n_25482, n_25483, n_25484, n_25485, n_25486, n_25487,
       n_25488;
  wire n_25489, n_25490, n_25491, n_25492, n_25493, n_25494, n_25495,
       n_25496;
  wire n_25497, n_25501, n_25502, n_25503, n_25504, n_25505, n_25506,
       n_25507;
  wire n_25508, n_25512, n_25513, n_25514, n_25515, n_25516, n_25517,
       n_25518;
  wire n_25519, n_25520, n_25521, n_25522, n_25523, n_25524, n_25525,
       n_25526;
  wire n_25527, n_25528, n_25529, n_25530, n_25531, n_25532, n_25533,
       n_25534;
  wire n_25543, n_25544, n_25545, n_25546, n_25547, n_25548, n_25549,
       n_25550;
  wire n_25551, n_25552, n_25553, n_25554, n_25555, n_25556, n_25557,
       n_25558;
  wire n_25559, n_25560, n_25561, n_25562, n_25563, n_25564, n_25565,
       n_25566;
  wire n_25567, n_25568, n_25569, n_25570, n_25571, n_25572, n_25573,
       n_25574;
  wire n_25575, n_25576, n_25577, n_25578, n_25579, n_25580, n_25581,
       n_25582;
  wire n_25583, n_25584, n_25585, n_25586, n_25587, n_25588, n_25589,
       n_25590;
  wire n_25591, n_25592, n_25593, n_25594, n_25595, n_25596, n_25597,
       n_25598;
  wire n_25599, n_25600, n_25601, n_25602, n_25603, n_25604, n_25605,
       n_25606;
  wire n_25607, n_25608, n_25609, n_25610, n_25611, n_25612, n_25613,
       n_25614;
  wire n_25615, n_25616, n_25617, n_25618, n_25619, n_25620, n_25621,
       n_25622;
  wire n_25623, n_25624, n_25625, n_25626, n_25627, n_25628, n_25629,
       n_25630;
  wire n_25631, n_25632, n_25633, n_25634, n_25635, n_25636, n_25637,
       n_25638;
  wire n_25639, n_25640, n_25641, n_25642, n_25643, n_25644, n_25645,
       n_25646;
  wire n_25647, n_25648, n_25649, n_25650, n_25651, n_25652, n_25653,
       n_25654;
  wire n_25655, n_25656, n_25657, n_25658, n_25659, n_25660, n_25661,
       n_25662;
  wire n_25663, n_25664, n_25665, n_25666, n_25667, n_25668, n_25669,
       n_25670;
  wire n_25671, n_25672, n_25673, n_25674, n_25675, n_25676, n_25677,
       n_25678;
  wire n_25679, n_25680, n_25681, n_25682, n_25683, n_25684, n_25685,
       n_25686;
  wire n_25687, n_25688, n_25689, n_25690, n_25691, n_25692, n_25693,
       n_25694;
  wire n_25695, n_25696, n_25697, n_25698, n_25699, n_25700, n_25701,
       n_25702;
  wire n_25703, n_25704, n_25705, n_25706, n_25707, n_25708, n_25709,
       n_25710;
  wire n_25711, n_25712, n_25713, n_25714, n_25715, n_25716, n_25717,
       n_25718;
  wire n_25719, n_25720, n_25721, n_25722, n_25723, n_25724, n_25725,
       n_25726;
  wire n_25727, n_25728, n_25729, n_25730, n_25731, n_25732, n_25733,
       n_25734;
  wire n_25735, n_25736, n_25737, n_25738, n_25739, n_25740, n_25741,
       n_25742;
  wire n_25743, n_25744, n_25745, n_25746, n_25747, n_25748, n_25749,
       n_25750;
  wire n_25751, n_25752, n_25753, n_25754, n_25755, n_25756, n_25757,
       n_25758;
  wire n_25759, n_25760, n_25761, n_25762, n_25763, n_25764, n_25765,
       n_25766;
  wire n_25767, n_25768, n_25769, n_25770, n_25771, n_25772, n_25773,
       n_25774;
  wire n_25775, n_25776, n_25777, n_25778, n_25779, n_25780, n_25781,
       n_25782;
  wire n_25783, n_25784, n_25785, n_25786, n_25787, n_25788, n_25789,
       n_25790;
  wire n_25791, n_25792, n_25793, n_25794, n_25795, n_25796, n_25797,
       n_25798;
  wire n_25799, n_25800, n_25801, n_25802, n_25803, n_25804, n_25805,
       n_25806;
  wire n_25807, n_25808, n_25809, n_25810, n_25811, n_25812, n_25813,
       n_25814;
  wire n_25815, n_25816, n_25817, n_25818, n_25819, n_25820, n_25821,
       n_25822;
  wire n_25823, n_25824, n_25825, n_25826, n_25827, n_25828, n_25829,
       n_25830;
  wire n_25831, n_25832, n_25833, n_25834, n_25835, n_25836, n_25837,
       n_25838;
  wire n_25839, n_25840, n_25841, n_25842, n_25843, n_25844, n_25845,
       n_25846;
  wire n_25847, n_25848, n_25849, n_25850, n_25851, n_25852, n_25853,
       n_25854;
  wire n_25855, n_25856, n_25857, n_25858, n_25859, n_25860, n_25861,
       n_25862;
  wire n_25863, n_25864, n_25865, n_25866, n_25867, n_25868, n_25869,
       n_25870;
  wire n_25871, n_25872, n_25873, n_25874, n_25875, n_25876, n_25877,
       n_25878;
  wire n_25879, n_25880, n_25881, n_25882, n_25883, n_25884, n_25885,
       n_25886;
  wire n_25887, n_25888, n_25889, n_25890, n_25891, n_25892, n_25893,
       n_25894;
  wire n_25895, n_25896, n_25897, n_25898, n_25899, n_25900, n_25901,
       n_25902;
  wire n_25903, n_25904, n_25905, n_25906, n_25907, n_25908, n_25909,
       n_25910;
  wire n_25911, n_25912, n_25913, n_25914, n_25915, n_25916, n_25917,
       n_25918;
  wire n_25919, n_25920, n_25921, n_25922, n_25923, n_25924, n_25925,
       n_25926;
  wire n_25927, n_25928, n_25929, n_25930, n_25931, n_25932, n_25933,
       n_25934;
  wire n_25935, n_25936, n_25937, n_25938, n_25939, n_25940, n_25941,
       n_25942;
  wire n_25943, n_25944, n_25945, n_25946, n_25947, n_25948, n_25949,
       n_25950;
  wire n_25951, n_25952, n_25953, n_25954, n_25955, n_25956, n_25957,
       n_25958;
  wire n_25959, n_25960, n_25961, n_25962, n_25963, n_25964, n_25965,
       n_25966;
  wire n_25967, n_25968, n_25969, n_25970, n_25971, n_25972, n_25973,
       n_25974;
  wire n_25975, n_25976, n_25977, n_25978, n_25979, n_25980, n_25981,
       n_25982;
  wire n_25983, n_25984, n_25985, n_25986, n_25987, n_25988, n_25989,
       n_25990;
  wire n_25991, n_25992, n_25993, n_25994, n_25995, n_25996, n_25997,
       n_25998;
  wire n_25999, n_26000, n_26001, n_26002, n_26003, n_26004, n_26005,
       n_26006;
  wire n_26007, n_26008, n_26009, n_26010, n_26011, n_26012, n_26013,
       n_26014;
  wire n_26015, n_26016, n_26017, n_26018, n_26019, n_26020, n_26021,
       n_26022;
  wire n_26023, n_26024, n_26025, n_26026, n_26027, n_26028, n_26029,
       n_26030;
  wire n_26031, n_26032, n_26033, n_26034, n_26035, n_26036, n_26037,
       n_26038;
  wire n_26039, n_26040, n_26041, n_26042, n_26043, n_26044, n_26045,
       n_26046;
  wire n_26047, n_26048, n_26049, n_26050, n_26051, n_26052, n_26053,
       n_26054;
  wire n_26055, n_26056, n_26057, n_26058, n_26059, n_26060, n_26061,
       n_26062;
  wire n_26063, n_26064, n_26065, n_26066, n_26067, n_26068, n_26069,
       n_26070;
  wire n_26071, n_26072, n_26073, n_26074, n_26075, n_26076, n_26077,
       n_26078;
  wire n_26079, n_26080, n_26081, n_26082, n_26083, n_26084, n_26085,
       n_26086;
  wire n_26087, n_26088, n_26089, n_26090, n_26091, n_26092, n_26093,
       n_26094;
  wire n_26095, n_26096, n_26097, n_26098, n_26099, n_26100, n_26101,
       n_26102;
  wire n_26103, n_26104, n_26105, n_26106, n_26107, n_26108, n_26109,
       n_26110;
  wire n_26111, n_26112, n_26113, n_26114, n_26115, n_26116, n_26117,
       n_26118;
  wire n_26119, n_26120, n_26121, n_26122, n_26123, n_26124, n_26125,
       n_26126;
  wire n_26127, n_26128, n_26129, n_26130, n_26131, n_26132, n_26133,
       n_26134;
  wire n_26135, n_26136, n_26137, n_26138, n_26139, n_26140, n_26141,
       n_26142;
  wire n_26143, n_26144, n_26145, n_26146, n_26147, n_26148, n_26149,
       n_26150;
  wire n_26151, n_26152, n_26153, n_26154, n_26155, n_26156, n_26158,
       n_26159;
  wire n_26160, n_26161, n_26162, n_26163, n_26164, n_26165, n_26166,
       n_26167;
  wire n_26168, n_26169, n_26170, n_26171, n_26172, n_26173, n_26174,
       n_26175;
  wire n_26176, n_26177, n_26178, n_26179, n_26180, n_26181, n_26182,
       n_26183;
  wire n_26184, n_26185, n_26186, n_26187, n_26188, n_26189, n_26190,
       n_26191;
  wire n_26192, n_26440, n_26441, n_26442, n_26443, n_26444, n_26445,
       n_26446;
  wire n_26447, n_26448, n_26449, n_26450, n_26451, n_26452, n_26453,
       n_26454;
  wire n_26455, n_26456, n_26457, n_26458, n_26459, n_26460, n_26461,
       n_26462;
  wire n_26463, n_26464, n_26465, n_26466, n_26467, n_26715, n_26716,
       n_26717;
  wire n_26718, n_26719, n_26720, n_26721, n_26722, n_26723, n_26724,
       n_26725;
  wire n_26726, n_26727, n_26728, n_26729, n_26730, n_26731, n_26732,
       n_26733;
  wire n_26734, n_26735, n_26736, n_26737, n_26738, n_26739, n_26740,
       n_26845;
  wire n_26846, n_26847, n_26848, n_26849, n_26850, n_26851, n_26852,
       n_26970;
  wire n_26971, n_26972, n_26973, n_26974, n_26975, n_26976, n_26977,
       n_26978;
  wire n_27096, n_27097, n_27098, n_27099, n_27100, n_27101, n_27102,
       n_27103;
  wire n_27104, n_27105, n_27106, n_27107, n_27108, n_27109, n_27110,
       n_27111;
  wire n_27112, n_27113, n_27114, n_27185, n_27186, n_27187, n_27188,
       n_27189;
  wire n_27190, n_27191, n_27192, n_27297, n_27298, n_27299, n_27300,
       n_27301;
  wire n_27302, n_27303, n_27304, n_27409, n_27410, n_27411, n_27412,
       n_27413;
  wire n_27414, n_27415, n_27416, n_27521, n_27522, n_27523, n_27524,
       n_27525;
  wire n_27526, n_27527, n_27528, n_27633, n_27634, n_27635, n_27636,
       n_27637;
  wire n_27638, n_27639, n_27640, n_27745, n_27746, n_27747, n_27748,
       n_27749;
  wire n_27750, n_27751, n_27752, n_27768, n_27769, n_27770, n_27771,
       n_27772;
  wire n_27773, n_27775, n_27776, n_27777, n_27779, n_27780, n_27781,
       n_27782;
  wire n_27785, n_27848, n_27852, n_27853, n_27859, n_27864, n_27870,
       n_27878;
  wire n_27879, n_27880, n_27882, n_27883, n_27963, n_27964, n_27967,
       n_27969;
  wire n_27977, n_27978, n_27981, n_27982, n_27983, n_27984, n_27985,
       n_27986;
  wire n_27991, n_27994, n_27995, n_27996, n_27997, n_27998, n_27999,
       n_28007;
  wire n_28008, n_28010, n_28011, n_28012, n_28014, n_28015, n_28017,
       n_28018;
  wire n_28019, n_28020, n_28021, n_28022, n_28023, n_28024, n_28025,
       n_28158;
  wire n_28159, n_28160, n_28161, n_28162, n_28163, n_28225, n_28226,
       n_28227;
  wire n_28228, n_28229, n_28230, n_28231, n_28232, n_28233, n_28234,
       n_28235;
  wire n_29266, n_29269, n_29270, n_29271, n_29272, n_29273, n_29274,
       n_29275;
  wire n_29276;
  fx68k_or_op g2(.A ({lineBmap[15], n_27782, n_27781, n_27780, n_27779,
       lineBmap[10], n_27777, n_27776, n_27775, 1'b0, n_27773, n_27772,
       n_27771, n_27770, n_27769, n_27768}), .Z (palIll));
  fx68k_or_op_4 g3(.A (opcode[7:0]), .Z (n_25805));
  fx68k_or_op_5 g4(.A (opcode[7:0]), .Z (n_25806));
  fx68k_case_box_16 ctl_178_19(.in_0 (col), .out_0 ({n_23482,
       UNCONNECTED3, n_23483, n_23484, n_23485, n_23486, n_23487,
       n_23488, n_23489, UNCONNECTED2, UNCONNECTED1, n_23490,
       UNCONNECTED0}));
  fx68k_mux_41 \mux_cmbsop_arA1[0]_178_19 (.ctl ({n_23482, n_23483,
       n_23484, n_23485, n_23486, n_23487, n_23488, n_23489, n_23490}),
       .in_0 (10'b0100000000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .in_8
       (10'b0111001100), .z ({\cmbsop_arA1[0] [19], \cmbsop_arA1[0]
       [18], \cmbsop_arA1[0] [17], \cmbsop_arA1[0] [16],
       \cmbsop_arA1[0] [15], \cmbsop_arA1[0] [14], \cmbsop_arA1[0]
       [13], \cmbsop_arA1[0] [12], \cmbsop_arA1[0] [11],
       \cmbsop_arA1[0] [10]}));
  fx68k_case_box_17 ctl_196_19(.in_0 (col), .out_0 ({n_23492,
       UNCONNECTED7, n_23493, n_23494, n_23495, n_23496, n_23497,
       n_23498, n_23499, UNCONNECTED6, UNCONNECTED5, n_23500,
       UNCONNECTED4}));
  fx68k_mux_41 \mux_cmbsop_arA1[0]_196_19 (.ctl ({n_23492, n_23493,
       n_23494, n_23495, n_23496, n_23497, n_23498, n_23499, n_23500}),
       .in_0 (10'b0100000000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .in_8
       (10'b0111001100), .z ({n_23954, n_23952, n_23950, n_23948,
       n_23946, n_23944, n_23942, n_23940, n_23938, n_23936}));
  fx68k_case_box_20 ctl_214_19(.in_0 (col), .out_0 ({n_23502,
       UNCONNECTED11, n_23503, n_23504, n_23505, n_23506, n_23507,
       n_23508, n_23509, UNCONNECTED10, UNCONNECTED9, n_23510,
       UNCONNECTED8}));
  fx68k_mux_41 \mux_cmbsop_arA1[0]_214_19 (.ctl ({n_23502, n_23503,
       n_23504, n_23505, n_23506, n_23507, n_23508, n_23509, n_23510}),
       .in_0 (10'b0100000000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .in_8
       (10'b0111001100), .z ({n_23934, n_23932, n_23930, n_23928,
       n_23926, n_23924, n_23922, n_23920, n_23918, n_23916}));
  fx68k_case_box_23 ctl_232_19(.in_0 (col), .out_0 ({n_23512,
       UNCONNECTED15, n_23513, n_23514, n_23515, n_23516, n_23517,
       n_23518, n_23519, UNCONNECTED14, UNCONNECTED13, n_23520,
       UNCONNECTED12}));
  fx68k_mux_41 \mux_cmbsop_arA1[0]_232_19 (.ctl ({n_23512, n_23513,
       n_23514, n_23515, n_23516, n_23517, n_23518, n_23519, n_23520}),
       .in_0 (10'b0100000000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .in_8
       (10'b0111001100), .z ({n_23914, n_23912, n_23910, n_23908,
       n_23906, n_23904, n_23902, n_23900, n_23898, n_23896}));
  fx68k_case_box_26 ctl_250_19(.in_0 (col), .out_0 ({n_23522,
       UNCONNECTED20, n_23523, n_23524, n_23525, n_23526, n_23527,
       n_23528, n_23529, UNCONNECTED19, UNCONNECTED18, UNCONNECTED17,
       UNCONNECTED16}));
  fx68k_mux_77 \mux_cmbsop_arA1[0]_250_19 (.ctl ({n_23522, n_23523,
       n_23524, n_23525, n_23526, n_23527, n_23528, n_23529}), .in_0
       (9'b100001100), .in_1 (9'b000001011), .in_2 (9'b000001111),
       .in_3 (9'b101111001), .in_4 (9'b111000110), .in_5
       (9'b111100111), .in_6 (9'b000001110), .in_7 (9'b111100110), .z
       ({n_23893, n_23891, n_23889, n_23887, n_23885, n_23883, n_23881,
       n_23879, n_23877}));
  fx68k_case_box_29 ctl_268_19(.in_0 (col), .out_0 ({n_23530,
       UNCONNECTED25, n_23531, n_23532, n_23533, n_23534, n_23535,
       n_23536, n_23537, UNCONNECTED24, UNCONNECTED23, UNCONNECTED22,
       UNCONNECTED21}));
  fx68k_mux_77 \mux_cmbsop_arA1[0]_268_19 (.ctl ({n_23530, n_23531,
       n_23532, n_23533, n_23534, n_23535, n_23536, n_23537}), .in_0
       (9'b100001100), .in_1 (9'b000001011), .in_2 (9'b000001111),
       .in_3 (9'b101111001), .in_4 (9'b111000110), .in_5
       (9'b111100111), .in_6 (9'b000001110), .in_7 (9'b111100110), .z
       ({n_23869, n_23864, n_23859, n_23854, n_23849, n_23844, n_23839,
       n_23834, n_23829}));
  fx68k_case_box_32 ctl_286_19(.in_0 (col), .out_0 ({n_23538,
       UNCONNECTED30, n_23539, n_23540, n_23541, n_23542, n_23543,
       n_23544, n_23545, UNCONNECTED29, UNCONNECTED28, UNCONNECTED27,
       UNCONNECTED26}));
  fx68k_mux_93 \mux_cmbsop_arA1[0]_286_19 (.ctl ({n_23538, n_23539,
       n_23540, n_23541, n_23542, n_23543, n_23544, n_23545}), .in_0
       (10'b0100000000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_23874, n_23870,
       n_23865, n_23860, n_23855, n_23850, n_23845, n_23840, n_23835,
       n_23830}));
  fx68k_case_box_35 ctl_304_19(.in_0 (col), .out_0 ({n_23546,
       UNCONNECTED35, n_23547, n_23548, n_23549, n_23550, n_23551,
       n_23552, n_23553, UNCONNECTED34, UNCONNECTED33, UNCONNECTED32,
       UNCONNECTED31}));
  fx68k_mux_93 \mux_cmbsop_arA1[0]_304_19 (.ctl ({n_23546, n_23547,
       n_23548, n_23549, n_23550, n_23551, n_23552, n_23553}), .in_0
       (10'b0100000000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_23875, n_23871,
       n_23866, n_23861, n_23856, n_23851, n_23846, n_23841, n_23836,
       n_23831}));
  fx68k_case_box_38 ctl_322_19(.in_0 (col), .out_0 ({n_23554,
       UNCONNECTED40, n_23555, n_23556, n_23557, n_23558, n_23559,
       n_23560, n_23561, UNCONNECTED39, UNCONNECTED38, UNCONNECTED37,
       UNCONNECTED36}));
  fx68k_mux_77 \mux_cmbsop_arA1[0]_322_19 (.ctl ({n_23554, n_23555,
       n_23556, n_23557, n_23558, n_23559, n_23560, n_23561}), .in_0
       (9'b100001100), .in_1 (9'b000001011), .in_2 (9'b000001111),
       .in_3 (9'b101111001), .in_4 (9'b111000110), .in_5
       (9'b111100111), .in_6 (9'b000001110), .in_7 (9'b111100110), .z
       ({n_23872, n_23867, n_23862, n_23857, n_23852, n_23847, n_23842,
       n_23837, n_23832}));
  fx68k_case_box_41 ctl_340_19(.in_0 (col), .out_0 ({n_23562, n_23563,
       n_23564, n_23565, n_23566, n_23567, n_23568, n_23569, n_23570,
       n_23571, n_23572, n_23573, UNCONNECTED41}));
  fx68k_mux_119 \mux_cmbsop_arA1[0]_340_19 (.ctl ({n_23562, n_23563,
       n_23564, n_23565, n_23566, n_23567, n_23568, n_23569, n_23570,
       n_23571, n_23572, n_23573}), .in_0 (10'b1111100111), .in_1
       (10'b0111010010), .in_2 (10'b0000000110), .in_3
       (10'b1000011100), .in_4 (10'b0100000011), .in_5
       (10'b0111000010), .in_6 (10'b0111100011), .in_7
       (10'b0000001010), .in_8 (10'b0111100010), .in_9
       (10'b0111000010), .in_10 (10'b0111100011), .in_11
       (10'b0011101010), .z ({n_25164, n_25159, n_25155, n_25150,
       n_25146, n_25141, n_25136, n_25132, n_25128, n_25123}));
  fx68k_case_box_44 ctl_358_19(.in_0 (col), .out_0 ({n_23574, n_23575,
       n_23576, n_23577, n_23578, n_23579, n_23580, n_23581, n_23582,
       UNCONNECTED45, UNCONNECTED44, UNCONNECTED43, UNCONNECTED42}));
  fx68k_mux_128 \mux_cmbsop_arA1[0]_358_19 (.ctl ({n_23574, n_23575,
       n_23576, n_23577, n_23578, n_23579, n_23580, n_23581, n_23582}),
       .in_0 (20'b11111011110000000000), .in_1
       (20'b01110101100000000000), .in_2 (20'b00000001100000000000),
       .in_3 (20'b10000111000000000000), .in_4
       (20'b01000000110000000000), .in_5 (20'b01110000100000000000),
       .in_6 (20'b01111000110000000000), .in_7
       (20'b00000010100000000000), .in_8 (20'b01111000100000000000), .z
       ({n_25165, n_25160, n_25156, n_25151, n_25147, n_25142, n_25137,
       n_25133, n_25129, n_25124, UNCONNECTED55, UNCONNECTED54,
       UNCONNECTED53, UNCONNECTED52, UNCONNECTED51, UNCONNECTED50,
       UNCONNECTED49, UNCONNECTED48, UNCONNECTED47, UNCONNECTED46}));
  fx68k_case_box_47 ctl_376_19(.in_0 (col), .out_0 ({n_23583, n_23584,
       n_23585, n_23586, n_23587, n_23588, n_23589, n_23590, n_23591,
       UNCONNECTED59, UNCONNECTED58, UNCONNECTED57, UNCONNECTED56}));
  fx68k_mux_128 \mux_cmbsop_arA1[0]_376_19 (.ctl ({n_23583, n_23584,
       n_23585, n_23586, n_23587, n_23588, n_23589, n_23590, n_23591}),
       .in_0 (20'b11111011110000000000), .in_1
       (20'b01110011100000000000), .in_2 (20'b00000001100000000000),
       .in_3 (20'b10000111000000000000), .in_4
       (20'b01000000110000000000), .in_5 (20'b01110000100000000000),
       .in_6 (20'b01111000110000000000), .in_7
       (20'b00000010100000000000), .in_8 (20'b01111000100000000000), .z
       ({n_25166, n_25161, n_25157, n_25152, n_25148, n_25143, n_25138,
       n_25134, n_25130, n_25125, UNCONNECTED69, UNCONNECTED68,
       UNCONNECTED67, UNCONNECTED66, UNCONNECTED65, UNCONNECTED64,
       UNCONNECTED63, UNCONNECTED62, UNCONNECTED61, UNCONNECTED60}));
  fx68k_case_box_50 ctl_394_19(.in_0 (col), .out_0 ({n_23592, n_23593,
       n_23594, n_23595, n_23596, n_23597, n_23598, n_23599, n_23600,
       UNCONNECTED73, UNCONNECTED72, UNCONNECTED71, UNCONNECTED70}));
  fx68k_mux_128 \mux_cmbsop_arA1[0]_394_19 (.ctl ({n_23592, n_23593,
       n_23594, n_23595, n_23596, n_23597, n_23598, n_23599, n_23600}),
       .in_0 (20'b11111010110000000000), .in_1
       (20'b01110010100000000000), .in_2 (20'b00000001100000000000),
       .in_3 (20'b10000111000000000000), .in_4
       (20'b01000000110000000000), .in_5 (20'b01110000100000000000),
       .in_6 (20'b01111000110000000000), .in_7
       (20'b00000010100000000000), .in_8 (20'b01111000100000000000), .z
       ({n_25167, n_25162, n_25158, n_25153, n_25149, n_25144, n_25139,
       n_25135, n_25131, n_25126, UNCONNECTED83, UNCONNECTED82,
       UNCONNECTED81, UNCONNECTED80, UNCONNECTED79, UNCONNECTED78,
       UNCONNECTED77, UNCONNECTED76, UNCONNECTED75, UNCONNECTED74}));
  fx68k_case_box_53 ctl_412_19(.in_0 (col), .out_0 ({n_23601,
       UNCONNECTED86, n_23602, n_23603, n_23604, n_23605, n_23606,
       n_23607, n_23608, n_23609, n_23610, UNCONNECTED85,
       UNCONNECTED84}));
  fx68k_mux_185 \mux_cmbsop_arA1[0]_412_19 (.ctl ({n_23601, n_23602,
       n_23603, n_23604, n_23605, n_23606, n_23607, n_23608, n_23609,
       n_23610}), .in_0 (10'b1111100111), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .in_8
       (10'b0111000010), .in_9 (10'b0111100011), .z ({n_23813, n_23806,
       n_23799, n_23792, n_23785, n_23778, n_23771, n_23764, n_23757,
       n_23750}));
  fx68k_case_box_56 ctl_430_19(.in_0 (col), .out_0 ({n_23611,
       UNCONNECTED91, n_23612, n_23613, n_23614, n_23615, n_23616,
       n_23617, n_23618, UNCONNECTED90, UNCONNECTED89, UNCONNECTED88,
       UNCONNECTED87}));
  fx68k_mux_93 \mux_cmbsop_arA1[0]_430_19 (.ctl ({n_23611, n_23612,
       n_23613, n_23614, n_23615, n_23616, n_23617, n_23618}), .in_0
       (10'b1111101111), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_23814, n_23807,
       n_23800, n_23793, n_23786, n_23779, n_23772, n_23765, n_23758,
       n_23751}));
  fx68k_case_box_59 ctl_448_19(.in_0 (col), .out_0 ({n_23619,
       UNCONNECTED96, n_23620, n_23621, n_23622, n_23623, n_23624,
       n_23625, n_23626, UNCONNECTED95, UNCONNECTED94, UNCONNECTED93,
       UNCONNECTED92}));
  fx68k_mux_93 \mux_cmbsop_arA1[0]_448_19 (.ctl ({n_23619, n_23620,
       n_23621, n_23622, n_23623, n_23624, n_23625, n_23626}), .in_0
       (10'b1111101111), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_23815, n_23808,
       n_23801, n_23794, n_23787, n_23780, n_23773, n_23766, n_23759,
       n_23752}));
  fx68k_case_box_62 ctl_466_19(.in_0 (col), .out_0 ({n_23627,
       UNCONNECTED101, n_23628, n_23629, n_23630, n_23631, n_23632,
       n_23633, n_23634, UNCONNECTED100, UNCONNECTED99, UNCONNECTED98,
       UNCONNECTED97}));
  fx68k_mux_93 \mux_cmbsop_arA1[0]_466_19 (.ctl ({n_23627, n_23628,
       n_23629, n_23630, n_23631, n_23632, n_23633, n_23634}), .in_0
       (10'b1111101011), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_23816, n_23809,
       n_23802, n_23795, n_23788, n_23781, n_23774, n_23767, n_23760,
       n_23753}));
  fx68k_case_box_65 ctl_484_19(.in_0 (col), .out_0 ({n_23635,
       UNCONNECTED106, n_23636, n_23637, n_23638, n_23639, n_23640,
       n_23641, n_23642, UNCONNECTED105, UNCONNECTED104,
       UNCONNECTED103, UNCONNECTED102}));
  fx68k_mux_93 \mux_cmbsop_arA1[0]_484_19 (.ctl ({n_23635, n_23636,
       n_23637, n_23638, n_23639, n_23640, n_23641, n_23642}), .in_0
       (10'b0100001000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_23817, n_23810,
       n_23803, n_23796, n_23789, n_23782, n_23775, n_23768, n_23761,
       n_23754}));
  fx68k_case_box_68 ctl_502_19(.in_0 (col), .out_0 ({n_23643,
       UNCONNECTED111, n_23644, n_23645, n_23646, n_23647, n_23648,
       n_23649, n_23650, UNCONNECTED110, UNCONNECTED109,
       UNCONNECTED108, UNCONNECTED107}));
  fx68k_mux_93 \mux_cmbsop_arA1[0]_502_19 (.ctl ({n_23643, n_23644,
       n_23645, n_23646, n_23647, n_23648, n_23649, n_23650}), .in_0
       (10'b0100001000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_23818, n_23811,
       n_23804, n_23797, n_23790, n_23783, n_23776, n_23769, n_23762,
       n_23755}));
  fx68k_case_box_71 ctl_520_19(.in_0 (col), .out_0 ({n_23651,
       UNCONNECTED116, n_23652, n_23653, n_23654, n_23655, n_23656,
       n_23657, n_23658, UNCONNECTED115, UNCONNECTED114,
       UNCONNECTED113, UNCONNECTED112}));
  fx68k_mux_77 \mux_cmbsop_arA1[0]_520_19 (.ctl ({n_23651, n_23652,
       n_23653, n_23654, n_23655, n_23656, n_23657, n_23658}), .in_0
       (9'b100000100), .in_1 (9'b000001011), .in_2 (9'b000001111),
       .in_3 (9'b101111001), .in_4 (9'b111000110), .in_5
       (9'b111100111), .in_6 (9'b000001110), .in_7 (9'b111100110), .z
       ({n_23812, n_23805, n_23798, n_23791, n_23784, n_23777, n_23770,
       n_23763, n_23756}));
  fx68k_mux_247 mux_scA3_411_10(.ctl ({n_23665, n_23666, n_23667,
       n_23668, n_23669, n_23670, n_23671}), .in_0 (8'b10001010), .in_1
       (8'b01000000), .in_2 (8'b01000000), .in_3 (8'b00110100), .in_4
       (8'b01000011), .in_5 (8'b01000011), .in_6 (8'b01000111), .z
       ({n_23690, n_23689, n_23688, n_23687, n_23686, n_23685, n_23684,
       n_23683}));
  fx68k_mux_254 mux_scA3_339_24(.ctl ({n_41, n_83, n_125, n_167,
       n_23682}), .in_0 (8'b10001010), .in_1 (8'b01000000), .in_2
       (8'b01000000), .in_3 (8'b00110100), .in_4 ({n_23690, n_23689,
       n_23688, n_23687, n_23686, n_23685, n_23684, n_23683}), .z
       ({n_23709, n_23708, n_23707, n_23706, n_23705, n_23704, n_23703,
       n_23702}));
  fx68k_mux_254 mux_scA3_267_24(.ctl ({n_23697, n_23698, n_23699,
       n_23700, n_23701}), .in_0 (8'b11001110), .in_1 (8'b11001100),
       .in_2 (8'b11001100), .in_3 (8'b11001110), .in_4 ({n_23709,
       n_23708, n_23707, n_23706, n_23705, n_23704, n_23703, n_23702}),
       .z ({n_23717, n_23716, n_23715, n_23714, n_23713, n_23712,
       n_23711, n_23710}));
  fx68k_bmux mux_scA3_249_32(.ctl (n_23521), .in_0 ({n_23717, n_23716,
       n_23715, n_23714, n_23713, n_23712, n_23711, n_23710}), .in_1
       (8'b11001110), .z ({n_23725, n_23724, n_23723, n_23722, n_23721,
       n_23720, n_23719, n_23718}));
  fx68k_bmux mux_scA3_231_32(.ctl (n_23511), .in_0 ({n_23725, n_23724,
       n_23723, n_23722, n_23721, n_23720, n_23719, n_23718}), .in_1
       (8'b11001100), .z ({n_23733, n_23732, n_23731, n_23730, n_23729,
       n_23728, n_23727, n_23726}));
  fx68k_bmux mux_scA3_213_32(.ctl (n_23501), .in_0 ({n_23733, n_23732,
       n_23731, n_23730, n_23729, n_23728, n_23727, n_23726}), .in_1
       (8'b11001100), .z ({n_23741, n_23740, n_23739, n_23738, n_23737,
       n_23736, n_23735, n_23734}));
  fx68k_bmux mux_scA3_195_32(.ctl (n_23491), .in_0 ({n_23741, n_23740,
       n_23739, n_23738, n_23737, n_23736, n_23735, n_23734}), .in_1
       (8'b11001100), .z ({n_23749, n_23748, n_23747, n_23746, n_23745,
       n_23744, n_23743, n_23742}));
  fx68k_bmux mux_scA3_177_27(.ctl (n_23477), .in_0 ({n_23749, n_23748,
       n_23747, n_23746, n_23745, n_23744, n_23743, n_23742}), .in_1
       (8'b11001100), .z ({scA3[9], scA3[7:1]}));
  fx68k_mux_272 \mux_arA23[0]_411_10 (.ctl ({n_23665, n_23666, n_23667,
       n_23668, n_23669, n_23670, n_23671}), .in_0 ({n_23813, n_23806,
       n_23799, n_23792, n_23785, n_23778, n_23771, n_23764, n_23757,
       n_23750}), .in_1 ({n_23814, n_23807, n_23800, n_23793, n_23786,
       n_23779, n_23772, n_23765, n_23758, n_23751}), .in_2 ({n_23815,
       n_23808, n_23801, n_23794, n_23787, n_23780, n_23773, n_23766,
       n_23759, n_23752}), .in_3 ({n_23816, n_23809, n_23802, n_23795,
       n_23788, n_23781, n_23774, n_23767, n_23760, n_23753}), .in_4
       ({n_23817, n_23810, n_23803, n_23796, n_23789, n_23782, n_23775,
       n_23768, n_23761, n_23754}), .in_5 ({n_23818, n_23811, n_23804,
       n_23797, n_23790, n_23783, n_23776, n_23769, n_23762, n_23755}),
       .in_6 ({1'b0, n_23812, n_23805, n_23798, n_23791, n_23784,
       n_23777, n_23770, n_23763, n_23756}), .z ({n_23828, n_23827,
       n_23826, n_23825, n_23824, n_23823, n_23822, n_23821, n_23820,
       n_23819}));
  fx68k_mux_281 \mux_arA23[0]_339_24 (.ctl ({n_41, n_23682}), .in_0
       (10'b0010101011), .in_1 ({n_23828, n_23827, n_23826, n_23825,
       n_23824, n_23823, n_23822, n_23821, n_23820, n_23819}), .z
       ({n_23876, n_23873, n_23868, n_23863, n_23858, n_23853, n_23848,
       n_23843, n_23838, n_23833}));
  fx68k_mux_290 \mux_arA23[0]_267_24 (.ctl ({n_23697, n_23698, n_23699,
       n_23700, n_23701}), .in_0 ({1'b0, n_23869, n_23864, n_23859,
       n_23854, n_23849, n_23844, n_23839, n_23834, n_23829}), .in_1
       ({n_23874, n_23870, n_23865, n_23860, n_23855, n_23850, n_23845,
       n_23840, n_23835, n_23830}), .in_2 ({n_23875, n_23871, n_23866,
       n_23861, n_23856, n_23851, n_23846, n_23841, n_23836, n_23831}),
       .in_3 ({1'b0, n_23872, n_23867, n_23862, n_23857, n_23852,
       n_23847, n_23842, n_23837, n_23832}), .in_4 ({n_23876, n_23873,
       n_23868, n_23863, n_23858, n_23853, n_23848, n_23843, n_23838,
       n_23833}), .z ({n_23895, n_23894, n_23892, n_23890, n_23888,
       n_23886, n_23884, n_23882, n_23880, n_23878}));
  fx68k_bmux_299 \mux_arA23[0]_249_32 (.ctl (n_23521), .in_0 ({n_23895,
       n_23894, n_23892, n_23890, n_23888, n_23886, n_23884, n_23882,
       n_23880, n_23878}), .in_1 ({1'b0, n_23893, n_23891, n_23889,
       n_23887, n_23885, n_23883, n_23881, n_23879, n_23877}), .z
       ({n_23915, n_23913, n_23911, n_23909, n_23907, n_23905, n_23903,
       n_23901, n_23899, n_23897}));
  fx68k_bmux_299 \mux_arA23[0]_231_32 (.ctl (n_23511), .in_0 ({n_23915,
       n_23913, n_23911, n_23909, n_23907, n_23905, n_23903, n_23901,
       n_23899, n_23897}), .in_1 ({n_23914, n_23912, n_23910, n_23908,
       n_23906, n_23904, n_23902, n_23900, n_23898, n_23896}), .z
       ({n_23935, n_23933, n_23931, n_23929, n_23927, n_23925, n_23923,
       n_23921, n_23919, n_23917}));
  fx68k_bmux_299 \mux_arA23[0]_213_32 (.ctl (n_23501), .in_0 ({n_23935,
       n_23933, n_23931, n_23929, n_23927, n_23925, n_23923, n_23921,
       n_23919, n_23917}), .in_1 ({n_23934, n_23932, n_23930, n_23928,
       n_23926, n_23924, n_23922, n_23920, n_23918, n_23916}), .z
       ({n_23955, n_23953, n_23951, n_23949, n_23947, n_23945, n_23943,
       n_23941, n_23939, n_23937}));
  fx68k_bmux_299 \mux_arA23[0]_195_32 (.ctl (n_23491), .in_0 ({n_23955,
       n_23953, n_23951, n_23949, n_23947, n_23945, n_23943, n_23941,
       n_23939, n_23937}), .in_1 ({n_23954, n_23952, n_23950, n_23948,
       n_23946, n_23944, n_23942, n_23940, n_23938, n_23936}), .z
       ({n_23965, n_23964, n_23963, n_23962, n_23961, n_23960, n_23959,
       n_23958, n_23957, n_23956}));
  fx68k_bmux_299 \mux_arA23[0]_177_27 (.ctl (n_23477), .in_0 ({n_23965,
       n_23964, n_23963, n_23962, n_23961, n_23960, n_23959, n_23958,
       n_23957, n_23956}), .in_1 ({\cmbsop_arA1[0] [19],
       \cmbsop_arA1[0] [18], \cmbsop_arA1[0] [17], \cmbsop_arA1[0]
       [16], \cmbsop_arA1[0] [15], \cmbsop_arA1[0] [14],
       \cmbsop_arA1[0] [13], \cmbsop_arA1[0] [12], \cmbsop_arA1[0]
       [11], \cmbsop_arA1[0] [10]}), .z ({\arA23[0] [9], \arA23[0] [8],
       \arA23[0] [7], \arA23[0] [6], \arA23[0] [5], \arA23[0] [4],
       \arA23[0] [3], \arA23[0] [2], \arA23[0] [1], \arA23[0] [0]}));
  fx68k_case_box_83 ctl_905_19(.in_0 (col), .out_0 ({n_23966,
       UNCONNECTED118, n_23967, n_23968, n_23969, n_23970, n_23971,
       n_23972, n_23973, n_23974, n_23975, n_23976, UNCONNECTED117}));
  fx68k_mux_304 \mux_cmbsop_arA1[1]_905_19 (.ctl ({n_23966, n_23967,
       n_23968, n_23969, n_23970, n_23971, n_23972, n_23973, n_23974,
       n_23975, n_23976}), .in_0 ({10'b0100100001, _X_, _X_, _X_, _X_,
       _X_, _X_, _X_}), .in_1 (17'b00000001101010111), .in_2
       (17'b10000111001010111), .in_3 (17'b01000000111010111), .in_4
       (17'b01110000101010111), .in_5 (17'b01111000111010111), .in_6
       (17'b00000010101010111), .in_7 (17'b01111000101010111), .in_8
       (17'b01110000101010111), .in_9 (17'b01111000111010111), .in_10
       (17'b00111010100101000), .z ({\cmbsop_arA1[1] [19],
       \cmbsop_arA1[1] [18], \cmbsop_arA1[1] [17], \cmbsop_arA1[1]
       [16], \cmbsop_arA1[1] [15], \cmbsop_arA1[1] [14],
       \cmbsop_arA1[1] [13], \cmbsop_arA1[1] [12], \cmbsop_arA1[1]
       [11], \cmbsop_arA1[1] [10], \cmbsop_arA1[1] [9],
       \cmbsop_arA1[1] [8], \cmbsop_arA1[1] [7], \cmbsop_arA1[1] [5],
       \cmbsop_arA1[1] [4], \cmbsop_arA1[1] [3], \cmbsop_arA1[1] [1]}));
  fx68k_case_box_86 ctl_922_19(.in_0 (col), .out_0 ({n_23977,
       UNCONNECTED120, n_23978, n_23979, n_23980, n_23981, n_23982,
       n_23983, n_23984, n_23985, n_23986, n_23987, UNCONNECTED119}));
  fx68k_mux_320 \mux_cmbsop_arA1[1]_922_19 (.ctl ({n_23977, n_23978,
       n_23979, n_23980, n_23981, n_23982, n_23983, n_23984, n_23985,
       n_23986, n_23987}), .in_0 ({10'b1011111010, _X_, _X_, _X_,
       _X_}), .in_1 (14'b00000001101001), .in_2 (14'b10000111001001),
       .in_3 (14'b01000000111001), .in_4 (14'b01110000101001), .in_5
       (14'b01111000111001), .in_6 (14'b00000010101001), .in_7
       (14'b01111000101001), .in_8 (14'b01110000101001), .in_9
       (14'b01111000111001), .in_10 (14'b00111010100110), .z ({n_25291,
       n_25284, n_25277, n_25270, n_25263, n_25256, n_25249, n_25242,
       n_25235, n_25228, n_24090, n_24082, n_24074, n_24066}));
  fx68k_case_box_89 ctl_939_19(.in_0 (col), .out_0 ({n_23988,
       UNCONNECTED122, n_23989, n_23990, n_23991, n_23992, n_23993,
       n_23994, n_23995, n_23996, n_23997, n_23998, UNCONNECTED121}));
  fx68k_mux_320 \mux_cmbsop_arA1[1]_939_19 (.ctl ({n_23988, n_23989,
       n_23990, n_23991, n_23992, n_23993, n_23994, n_23995, n_23996,
       n_23997, n_23998}), .in_0 ({10'b1011111110, _X_, _X_, _X_,
       _X_}), .in_1 (14'b00000001101001), .in_2 (14'b10000111001001),
       .in_3 (14'b01000000111001), .in_4 (14'b01110000101001), .in_5
       (14'b01111000111001), .in_6 (14'b00000010101001), .in_7
       (14'b01111000101001), .in_8 (14'b01110000101001), .in_9
       (14'b01111000111001), .in_10 (14'b00111010100110), .z ({n_25292,
       n_25285, n_25278, n_25271, n_25264, n_25257, n_25250, n_25243,
       n_25236, n_25229, n_24091, n_24083, n_24075, n_24067}));
  fx68k_case_box_92 ctl_956_19(.in_0 (col), .out_0 ({n_23999,
       UNCONNECTED124, n_24000, n_24001, n_24002, n_24003, n_24004,
       n_24005, n_24006, n_24007, n_24008, n_24009, UNCONNECTED123}));
  fx68k_mux_346 \mux_cmbsop_arA1[1]_956_19 (.ctl ({n_23999, n_24000,
       n_24001, n_24002, n_24003, n_24004, n_24005, n_24006, n_24007,
       n_24008, n_24009}), .in_0 ({10'b1011111000, _X_, _X_, _X_, _X_,
       _X_, _X_}), .in_1 (16'b0000000110100011), .in_2
       (16'b1000011100100011), .in_3 (16'b0100000011100011), .in_4
       (16'b0111000010100011), .in_5 (16'b0111100011100011), .in_6
       (16'b0000001010100011), .in_7 (16'b0111100010100011), .in_8
       (16'b0111000010100011), .in_9 (16'b0111100011100011), .in_10
       (16'b0011101010011100), .z ({n_25293, n_25286, n_25279, n_25272,
       n_25265, n_25258, n_25251, n_25244, n_25237, n_25230, n_24092,
       n_24084, n_24080, n_24076, n_24072, n_24068}));
  fx68k_case_box_95 ctl_973_19(.in_0 (col), .out_0 ({n_24010,
       UNCONNECTED126, n_24011, n_24012, n_24013, n_24014, n_24015,
       n_24016, n_24017, n_24018, n_24019, n_24020, UNCONNECTED125}));
  fx68k_mux_361 \mux_cmbsop_arA1[1]_973_19 (.ctl ({n_24010, n_24011,
       n_24012, n_24013, n_24014, n_24015, n_24016, n_24017, n_24018,
       n_24019, n_24020}), .in_0 ({10'b1011011010, _X_, _X_, _X_}),
       .in_1 (13'b0000000110100), .in_2 (13'b1000011100100), .in_3
       (13'b0100000011100), .in_4 (13'b0111000010100), .in_5
       (13'b0111100011100), .in_6 (13'b0000001010100), .in_7
       (13'b0111100010100), .in_8 (13'b0111000010100), .in_9
       (13'b0111100011100), .in_10 (13'b0011101010011), .z ({n_25294,
       n_25287, n_25280, n_25273, n_25266, n_25259, n_25252, n_25245,
       n_25238, n_25231, n_24093, n_24085, n_24077}));
  fx68k_case_box_98 ctl_990_19(.in_0 (col), .out_0 ({n_24021,
       UNCONNECTED128, n_24022, n_24023, n_24024, n_24025, n_24026,
       n_24027, n_24028, n_24029, n_24030, n_24031, UNCONNECTED127}));
  fx68k_mux_304 \mux_cmbsop_arA1[1]_990_19 (.ctl ({n_24021, n_24022,
       n_24023, n_24024, n_24025, n_24026, n_24027, n_24028, n_24029,
       n_24030, n_24031}), .in_0 ({10'b0111101011, _X_, _X_, _X_, _X_,
       _X_, _X_, _X_}), .in_1 (17'b00000001101000100), .in_2
       (17'b10000111001000100), .in_3 (17'b01000000111000100), .in_4
       (17'b01110000101000100), .in_5 (17'b01111000111000100), .in_6
       (17'b00000010101000100), .in_7 (17'b01111000101000100), .in_8
       (17'b01110000101000100), .in_9 (17'b01111000111000100), .in_10
       (17'b00111010100111011), .z ({n_25295, n_25288, n_25281,
       n_25274, n_25267, n_25260, n_25253, n_25246, n_25239, n_25232,
       n_24096, n_24094, n_24086, n_24081, n_24078, n_24073, n_24069}));
  fx68k_case_box_101 ctl_1007_19(.in_0 (col), .out_0 ({n_24032,
       UNCONNECTED130, n_24033, n_24034, n_24035, n_24036, n_24037,
       n_24038, n_24039, n_24040, n_24041, n_24042, UNCONNECTED129}));
  fx68k_mux_320 \mux_cmbsop_arA1[1]_1007_19 (.ctl ({n_24032, n_24033,
       n_24034, n_24035, n_24036, n_24037, n_24038, n_24039, n_24040,
       n_24041, n_24042}), .in_0 ({10'b1011011001, _X_, _X_, _X_,
       _X_}), .in_1 (14'b00000001101000), .in_2 (14'b10000111001000),
       .in_3 (14'b01000000111000), .in_4 (14'b01110000101000), .in_5
       (14'b01111000111000), .in_6 (14'b00000010101000), .in_7
       (14'b01111000101000), .in_8 (14'b01110000101000), .in_9
       (14'b01111000111000), .in_10 (14'b00111010100111), .z ({n_25296,
       n_25289, n_25282, n_25275, n_25268, n_25261, n_25254, n_25247,
       n_25240, n_25233, n_24095, n_24087, n_24079, n_24070}));
  fx68k_case_box_104 ctl_1024_19(.in_0 (col), .out_0 ({n_24043,
       UNCONNECTED132, n_24044, n_24045, n_24046, n_24047, n_24048,
       n_24049, n_24050, n_24051, n_24052, n_24053, UNCONNECTED131}));
  fx68k_mux_320 \mux_cmbsop_arA1[1]_1024_19 (.ctl ({n_24043, n_24044,
       n_24045, n_24046, n_24047, n_24048, n_24049, n_24050, n_24051,
       n_24052, n_24053}), .in_0 ({10'b0111101010, _X_, _X_, _X_,
       _X_}), .in_1 (14'b00000001101001), .in_2 (14'b10000111001001),
       .in_3 (14'b01000000111001), .in_4 (14'b01110000101001), .in_5
       (14'b01111000111001), .in_6 (14'b00000010101001), .in_7
       (14'b01111000101001), .in_8 (14'b01110000101001), .in_9
       (14'b01111000111001), .in_10 (14'b00111010100110), .z ({n_25297,
       n_25290, n_25283, n_25276, n_25269, n_25262, n_25255, n_25248,
       n_25241, n_25234, n_24097, n_24089, n_24088, n_24071}));
  fx68k_mux_93 \mux_arA23[1]_902_14 (.ctl ({n_24058, n_24059, n_24060,
       n_24061, n_24062, n_24063, n_24064, n_24065}), .in_0
       ({\cmbsop_arA1[1] [9], \cmbsop_arA1[1] [8], \cmbsop_arA1[1] [7],
       1'b0, \cmbsop_arA1[1] [5], \cmbsop_arA1[1] [4],
       \cmbsop_arA1[1] [3], 1'b0, \cmbsop_arA1[1] [1], 1'b1}), .in_1
       ({1'b1, n_24090, 1'b1, n_24082, 1'b1, n_24074, 3'b101,
       n_24066}), .in_2 ({1'b1, n_24091, 1'b1, n_24083, 1'b1, n_24075,
       3'b111, n_24067}), .in_3 ({1'b1, n_24092, 1'b1, n_24084,
       n_24080, n_24076, 2'b10, n_24072, n_24068}), .in_4 ({1'b1,
       n_24093, 1'b1, n_24085, 1'b0, n_24077, 4'b1010}), .in_5
       ({n_24096, n_24094, 1'b1, n_24086, n_24081, n_24078, 2'b10,
       n_24073, n_24069}), .in_6 ({1'b1, n_24095, 1'b1, n_24087, 1'b0,
       n_24079, 3'b100, n_24070}), .in_7 ({n_24097, 1'b1, n_24089,
       n_24088, 5'b10101, n_24071}), .z ({\arA23[1] [9], \arA23[1] [8],
       \arA23[1] [7], \arA23[1] [6], \arA23[1] [5], \arA23[1] [4],
       \arA23[1] [3], \arA23[1] [2], \arA23[1] [1], \arA23[1] [0]}));
  fx68k_case_box_110 ctl_1048_19(.in_0 (col), .out_0 ({n_24098,
       n_24099, n_24100, n_24101, n_24102, n_24103, n_24104, n_24105,
       n_24106, n_24107, n_24108, n_24109, UNCONNECTED133}));
  fx68k_mux_424 \mux_cmbsop_arA1[2]_1048_19 (.ctl ({n_24098, n_24099,
       n_24100, n_24101, n_24102, n_24103, n_24104, n_24105, n_24106,
       n_24107, n_24108, n_24109}), .in_0 ({9'b100101001, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_1 ({9'b100101001, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_2 (16'b0000010111010111), .in_3
       (16'b0000011111010111), .in_4 (16'b1011110011010111), .in_5
       (16'b1110001101010111), .in_6 (16'b1111001111010111), .in_7
       (16'b0000011101010111), .in_8 (16'b1111001101010111), .in_9
       (16'b1110001101010111), .in_10 (16'b1111001111010111), .in_11
       (16'b0101001110101000), .z ({\cmbsop_arA1[2] [18],
       \cmbsop_arA1[2] [17], \cmbsop_arA1[2] [16], \cmbsop_arA1[2]
       [15], \cmbsop_arA1[2] [14], \cmbsop_arA1[2] [13],
       \cmbsop_arA1[2] [12], \cmbsop_arA1[2] [11], \cmbsop_arA1[2]
       [10], \cmbsop_arA1[2] [9], \cmbsop_arA1[2] [8],
       \cmbsop_arA1[2] [7], \cmbsop_arA1[2] [5], \cmbsop_arA1[2] [4],
       \cmbsop_arA1[2] [2], \cmbsop_arA1[2] [1]}));
  fx68k_case_box_113 ctl_1065_19(.in_0 (col), .out_0 ({n_24110,
       n_24111, n_24112, n_24113, n_24114, n_24115, n_24116, n_24117,
       n_24118, n_24119, n_24120, n_24121, UNCONNECTED134}));
  fx68k_mux_424 \mux_cmbsop_arA1[2]_1065_19 (.ctl ({n_24110, n_24111,
       n_24112, n_24113, n_24114, n_24115, n_24116, n_24117, n_24118,
       n_24119, n_24120, n_24121}), .in_0 ({9'b100101001, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_1 ({9'b100101001, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_2 (16'b0000010111010111), .in_3
       (16'b0000011111010111), .in_4 (16'b1011110011010111), .in_5
       (16'b1110001101010111), .in_6 (16'b1111001111010111), .in_7
       (16'b0000011101010111), .in_8 (16'b1111001101010111), .in_9
       (16'b1110001101010111), .in_10 (16'b1111001111010111), .in_11
       (16'b0101001110101000), .z ({n_25362, n_25354, n_25346, n_25338,
       n_25330, n_25322, n_25314, n_25306, n_25298, n_24241, n_24234,
       n_24232, n_24221, n_24214, n_24213, n_24210}));
  fx68k_case_box_116 ctl_1082_19(.in_0 (col), .out_0 ({n_24122,
       n_24123, n_24124, n_24125, n_24126, n_24127, n_24128, n_24129,
       n_24130, n_24131, n_24132, n_24133, UNCONNECTED135}));
  fx68k_mux_454 \mux_cmbsop_arA1[2]_1082_19 (.ctl ({n_24122, n_24123,
       n_24124, n_24125, n_24126, n_24127, n_24128, n_24129, n_24130,
       n_24131, n_24132, n_24133}), .in_0 ({10'b1011111001, _X_, _X_,
       _X_}), .in_1 ({10'b1011111001, _X_, _X_, _X_}), .in_2
       (13'b0000001011100), .in_3 (13'b0000001111100), .in_4
       (13'b0101111001100), .in_5 (13'b0111000110100), .in_6
       (13'b0111100111100), .in_7 (13'b0000001110100), .in_8
       (13'b0111100110100), .in_9 (13'b0111000110100), .in_10
       (13'b0111100111100), .in_11 (13'b0010100111011), .z ({n_25370,
       n_25363, n_25355, n_25347, n_25339, n_25331, n_25323, n_25315,
       n_25307, n_25299, n_24235, n_24225, n_24215}));
  fx68k_case_box_119 ctl_1099_19(.in_0 (col), .out_0 ({n_24134,
       n_24135, n_24136, n_24137, n_24138, n_24139, n_24140, n_24141,
       n_24142, n_24143, n_24144, n_24145, UNCONNECTED136}));
  fx68k_mux_454 \mux_cmbsop_arA1[2]_1099_19 (.ctl ({n_24134, n_24135,
       n_24136, n_24137, n_24138, n_24139, n_24140, n_24141, n_24142,
       n_24143, n_24144, n_24145}), .in_0 ({10'b1011111101, _X_, _X_,
       _X_}), .in_1 ({10'b1011111101, _X_, _X_, _X_}), .in_2
       (13'b0000001011100), .in_3 (13'b0000001111100), .in_4
       (13'b0101111001100), .in_5 (13'b0111000110100), .in_6
       (13'b0111100111100), .in_7 (13'b0000001110100), .in_8
       (13'b0111100110100), .in_9 (13'b0111000110100), .in_10
       (13'b0111100111100), .in_11 (13'b0010100111011), .z ({n_25371,
       n_25364, n_25356, n_25348, n_25340, n_25332, n_25324, n_25316,
       n_25308, n_25300, n_24236, n_24226, n_24216}));
  fx68k_case_box_122 ctl_1116_19(.in_0 (col), .out_0 ({n_24146,
       n_24147, n_24148, n_24149, n_24150, n_24151, n_24152, n_24153,
       n_24154, n_24155, n_24156, n_24157, UNCONNECTED137}));
  fx68k_mux_424 \mux_cmbsop_arA1[2]_1116_19 (.ctl ({n_24146, n_24147,
       n_24148, n_24149, n_24150, n_24151, n_24152, n_24153, n_24154,
       n_24155, n_24156, n_24157}), .in_0 ({10'b1011111100, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_1 ({10'b1011111100, _X_, _X_, _X_,
       _X_, _X_, _X_}), .in_2 (16'b0000001011100011), .in_3
       (16'b0000001111100011), .in_4 (16'b0101111001100011), .in_5
       (16'b0111000110100011), .in_6 (16'b0111100111100011), .in_7
       (16'b0000001110100011), .in_8 (16'b0111100110100011), .in_9
       (16'b0111000110100011), .in_10 (16'b0111100111100011), .in_11
       (16'b0010100111011100), .z ({n_25372, n_25365, n_25357, n_25349,
       n_25341, n_25333, n_25325, n_25317, n_25309, n_25301, n_24237,
       n_24227, n_24222, n_24217, n_24211, n_24206}));
  fx68k_case_box_125 ctl_1133_19(.in_0 (col), .out_0 ({n_24158,
       n_24159, n_24160, n_24161, n_24162, n_24163, n_24164, n_24165,
       n_24166, n_24167, n_24168, n_24169, UNCONNECTED138}));
  fx68k_mux_454 \mux_cmbsop_arA1[2]_1133_19 (.ctl ({n_24158, n_24159,
       n_24160, n_24161, n_24162, n_24163, n_24164, n_24165, n_24166,
       n_24167, n_24168, n_24169}), .in_0 ({10'b1011011110, _X_, _X_,
       _X_}), .in_1 ({10'b1011011110, _X_, _X_, _X_}), .in_2
       (13'b0000001011100), .in_3 (13'b0000001111100), .in_4
       (13'b0101111001100), .in_5 (13'b0111000110100), .in_6
       (13'b0111100111100), .in_7 (13'b0000001110100), .in_8
       (13'b0111100110100), .in_9 (13'b0111000110100), .in_10
       (13'b0111100111100), .in_11 (13'b0010100111011), .z ({n_25373,
       n_25366, n_25358, n_25350, n_25342, n_25334, n_25326, n_25318,
       n_25310, n_25302, n_24238, n_24228, n_24218}));
  fx68k_case_box_128 ctl_1150_19(.in_0 (col), .out_0 ({n_24170,
       n_24171, n_24172, n_24173, n_24174, n_24175, n_24176, n_24177,
       n_24178, n_24179, n_24180, n_24181, UNCONNECTED139}));
  fx68k_mux_424 \mux_cmbsop_arA1[2]_1150_19 (.ctl ({n_24170, n_24171,
       n_24172, n_24173, n_24174, n_24175, n_24176, n_24177, n_24178,
       n_24179, n_24180, n_24181}), .in_0 ({9'b111101111, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_1 ({9'b111101111, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_2 (16'b0000010111000100), .in_3
       (16'b0000011111000100), .in_4 (16'b1011110011000100), .in_5
       (16'b1110001101000100), .in_6 (16'b1111001111000100), .in_7
       (16'b0000011101000100), .in_8 (16'b1111001101000100), .in_9
       (16'b1110001101000100), .in_10 (16'b1111001111000100), .in_11
       (16'b0101001110111011), .z ({n_25367, n_25359, n_25351, n_25343,
       n_25335, n_25327, n_25319, n_25311, n_25303, n_24242, n_24239,
       n_24229, n_24223, n_24219, n_24212, n_24207}));
  fx68k_case_box_131 ctl_1167_19(.in_0 (col), .out_0 ({n_24182,
       n_24183, n_24184, n_24185, n_24186, n_24187, n_24188, n_24189,
       n_24190, n_24191, n_24192, n_24193, UNCONNECTED140}));
  fx68k_mux_520 \mux_cmbsop_arA1[2]_1167_19 (.ctl ({n_24182, n_24183,
       n_24184, n_24185, n_24186, n_24187, n_24188, n_24189, n_24190,
       n_24191, n_24192, n_24193}), .in_0 ({10'b1011011101, _X_, _X_,
       _X_, _X_}), .in_1 ({10'b1011011101, _X_, _X_, _X_, _X_}), .in_2
       (14'b00000010111000), .in_3 (14'b00000011111000), .in_4
       (14'b01011110011000), .in_5 (14'b01110001101000), .in_6
       (14'b01111001111000), .in_7 (14'b00000011101000), .in_8
       (14'b01111001101000), .in_9 (14'b01110001101000), .in_10
       (14'b01111001111000), .in_11 (14'b00101001110111), .z ({n_25374,
       n_25368, n_25360, n_25352, n_25344, n_25336, n_25328, n_25320,
       n_25312, n_25304, n_24240, n_24230, n_24220, n_24208}));
  fx68k_case_box_134 ctl_1184_19(.in_0 (col), .out_0 ({n_24194,
       n_24195, n_24196, n_24197, n_24198, n_24199, n_24200, n_24201,
       n_24202, n_24203, n_24204, n_24205, UNCONNECTED141}));
  fx68k_mux_520 \mux_cmbsop_arA1[2]_1184_19 (.ctl ({n_24194, n_24195,
       n_24196, n_24197, n_24198, n_24199, n_24200, n_24201, n_24202,
       n_24203, n_24204, n_24205}), .in_0 ({9'b111101110, _X_, _X_,
       _X_, _X_, _X_}), .in_1 ({9'b111101110, _X_, _X_, _X_, _X_,
       _X_}), .in_2 (14'b00000101110001), .in_3 (14'b00000111110001),
       .in_4 (14'b10111100110001), .in_5 (14'b11100011010001), .in_6
       (14'b11110011110001), .in_7 (14'b00000111010001), .in_8
       (14'b11110011010001), .in_9 (14'b11100011010001), .in_10
       (14'b11110011110001), .in_11 (14'b01010011101110), .z ({n_25369,
       n_25361, n_25353, n_25345, n_25337, n_25329, n_25321, n_25313,
       n_25305, n_24243, n_24233, n_24231, n_24224, n_24209}));
  fx68k_bmux_546 \mux_arA23[2]_1045_14 (.ctl (movEa), .in_0
       ({\cmbsop_arA1[2] [9], \cmbsop_arA1[2] [8], \cmbsop_arA1[2] [7],
       1'b0, \cmbsop_arA1[2] [5], \cmbsop_arA1[2] [4],
       \cmbsop_arA1[2] [2], \cmbsop_arA1[2] [1], 1'b1}), .in_1
       ({n_24241, n_24234, n_24232, 1'b0, n_24221, n_24214, n_24213,
       n_24210, 1'b1}), .in_2 ({1'b1, n_24235, 1'b1, n_24225, 1'b1,
       n_24215, 3'b001}), .in_3 ({1'b1, n_24236, 1'b1, n_24226, 1'b1,
       n_24216, 3'b101}), .in_4 ({1'b1, n_24237, 1'b1, n_24227,
       n_24222, n_24217, 1'b1, n_24211, n_24206}), .in_5 ({1'b1,
       n_24238, 1'b1, n_24228, 1'b0, n_24218, 3'b110}), .in_6
       ({n_24242, n_24239, 1'b1, n_24229, n_24223, n_24219, 1'b1,
       n_24212, n_24207}), .in_7 ({1'b1, n_24240, 1'b1, n_24230, 1'b0,
       n_24220, 2'b10, n_24208}), .in_8 ({n_24243, 1'b1, n_24233,
       n_24231, n_24224, 3'b011, n_24209}), .z ({\arA23[2] [9],
       \arA23[2] [8], \arA23[2] [7], \arA23[2] [6], \arA23[2] [5],
       \arA23[2] [4], \arA23[2] [2], \arA23[2] [1], \arA23[2] [0]}));
  fx68k_case_box_137 ctl_1208_19(.in_0 (col), .out_0 ({n_24244,
       n_24245, n_24246, n_24247, n_24248, n_24249, n_24250, n_24251,
       n_24252, n_24253, n_24254, n_24255, UNCONNECTED142}));
  fx68k_mux_547 \mux_cmbsop_arA1[3]_1208_19 (.ctl ({n_24244, n_24245,
       n_24246, n_24247, n_24248, n_24249, n_24250, n_24251, n_24252,
       n_24253, n_24254, n_24255}), .in_0 ({10'b0100100001, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_1 ({10'b0100100001, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_2 (17'b00000001101010111), .in_3
       (17'b10000111001010111), .in_4 (17'b01000000111010111), .in_5
       (17'b01110000101010111), .in_6 (17'b01111000111010111), .in_7
       (17'b00000010101010111), .in_8 (17'b01111000101010111), .in_9
       (17'b01110000101010111), .in_10 (17'b01111000111010111), .in_11
       (17'b00111010100101000), .z ({\cmbsop_arA1[3] [19],
       \cmbsop_arA1[3] [18], \cmbsop_arA1[3] [17], \cmbsop_arA1[3]
       [16], \cmbsop_arA1[3] [15], \cmbsop_arA1[3] [14],
       \cmbsop_arA1[3] [13], \cmbsop_arA1[3] [12], \cmbsop_arA1[3]
       [11], \cmbsop_arA1[3] [10], \cmbsop_arA1[3] [9],
       \cmbsop_arA1[3] [8], \cmbsop_arA1[3] [7], \cmbsop_arA1[3] [5],
       \cmbsop_arA1[3] [4], \cmbsop_arA1[3] [3], \cmbsop_arA1[3] [1]}));
  fx68k_case_box_140 ctl_1225_19(.in_0 (col), .out_0 ({n_24256,
       n_24257, n_24258, n_24259, n_24260, n_24261, n_24262, n_24263,
       n_24264, n_24265, n_24266, n_24267, UNCONNECTED143}));
  fx68k_mux_520 \mux_cmbsop_arA1[3]_1225_19 (.ctl ({n_24256, n_24257,
       n_24258, n_24259, n_24260, n_24261, n_24262, n_24263, n_24264,
       n_24265, n_24266, n_24267}), .in_0 ({10'b1001111001, _X_, _X_,
       _X_, _X_}), .in_1 ({10'b1001111001, _X_, _X_, _X_, _X_}), .in_2
       (14'b00000001100100), .in_3 (14'b10000111000100), .in_4
       (14'b01000000110100), .in_5 (14'b01110000100100), .in_6
       (14'b01111000110100), .in_7 (14'b00000010100100), .in_8
       (14'b01111000100100), .in_9 (14'b01110000100100), .in_10
       (14'b01111000110100), .in_11 (14'b00111010101011), .z ({n_25447,
       n_25439, n_25431, n_25423, n_25415, n_25407, n_25399, n_25391,
       n_25383, n_25375, n_24394, n_24387, n_24376, n_24361}));
  fx68k_case_box_143 ctl_1242_19(.in_0 (col), .out_0 ({n_24268,
       n_24269, n_24270, n_24271, n_24272, n_24273, n_24274, n_24275,
       n_24276, n_24277, n_24278, n_24279, UNCONNECTED144}));
  fx68k_mux_520 \mux_cmbsop_arA1[3]_1242_19 (.ctl ({n_24268, n_24269,
       n_24270, n_24271, n_24272, n_24273, n_24274, n_24275, n_24276,
       n_24277, n_24278, n_24279}), .in_0 ({10'b1011111010, _X_, _X_,
       _X_, _X_}), .in_1 ({10'b1011111010, _X_, _X_, _X_, _X_}), .in_2
       (14'b00000001101001), .in_3 (14'b10000111001001), .in_4
       (14'b01000000111001), .in_5 (14'b01110000101001), .in_6
       (14'b01111000111001), .in_7 (14'b00000010101001), .in_8
       (14'b01111000101001), .in_9 (14'b01110000101001), .in_10
       (14'b01111000111001), .in_11 (14'b00111010100110), .z ({n_25448,
       n_25440, n_25432, n_25424, n_25416, n_25408, n_25400, n_25392,
       n_25384, n_25376, n_24388, n_24379, n_24370, n_24362}));
  fx68k_case_box_146 ctl_1259_19(.in_0 (col), .out_0 ({n_24280,
       n_24281, n_24282, n_24283, n_24284, n_24285, n_24286, n_24287,
       n_24288, n_24289, n_24290, n_24291, UNCONNECTED145}));
  fx68k_mux_520 \mux_cmbsop_arA1[3]_1259_19 (.ctl ({n_24280, n_24281,
       n_24282, n_24283, n_24284, n_24285, n_24286, n_24287, n_24288,
       n_24289, n_24290, n_24291}), .in_0 ({10'b1011111110, _X_, _X_,
       _X_, _X_}), .in_1 ({10'b1011111110, _X_, _X_, _X_, _X_}), .in_2
       (14'b00000001101001), .in_3 (14'b10000111001001), .in_4
       (14'b01000000111001), .in_5 (14'b01110000101001), .in_6
       (14'b01111000111001), .in_7 (14'b00000010101001), .in_8
       (14'b01111000101001), .in_9 (14'b01110000101001), .in_10
       (14'b01111000111001), .in_11 (14'b00111010100110), .z ({n_25449,
       n_25441, n_25433, n_25425, n_25417, n_25409, n_25401, n_25393,
       n_25385, n_25377, n_24389, n_24380, n_24371, n_24363}));
  fx68k_case_box_149 ctl_1276_19(.in_0 (col), .out_0 ({n_24292,
       n_24293, n_24294, n_24295, n_24296, n_24297, n_24298, n_24299,
       n_24300, n_24301, n_24302, n_24303, UNCONNECTED146}));
  fx68k_mux_424 \mux_cmbsop_arA1[3]_1276_19 (.ctl ({n_24292, n_24293,
       n_24294, n_24295, n_24296, n_24297, n_24298, n_24299, n_24300,
       n_24301, n_24302, n_24303}), .in_0 ({10'b1011111000, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_1 ({10'b1011111000, _X_, _X_, _X_,
       _X_, _X_, _X_}), .in_2 (16'b0000000110100011), .in_3
       (16'b1000011100100011), .in_4 (16'b0100000011100011), .in_5
       (16'b0111000010100011), .in_6 (16'b0111100011100011), .in_7
       (16'b0000001010100011), .in_8 (16'b0111100010100011), .in_9
       (16'b0111000010100011), .in_10 (16'b0111100011100011), .in_11
       (16'b0011101010011100), .z ({n_25450, n_25442, n_25434, n_25426,
       n_25418, n_25410, n_25402, n_25394, n_25386, n_25378, n_24390,
       n_24381, n_24377, n_24372, n_24368, n_24364}));
  fx68k_case_box_152 ctl_1293_19(.in_0 (col), .out_0 ({n_24304,
       n_24305, n_24306, n_24307, n_24308, n_24309, n_24310, n_24311,
       n_24312, n_24313, n_24314, n_24315, UNCONNECTED147}));
  fx68k_mux_454 \mux_cmbsop_arA1[3]_1293_19 (.ctl ({n_24304, n_24305,
       n_24306, n_24307, n_24308, n_24309, n_24310, n_24311, n_24312,
       n_24313, n_24314, n_24315}), .in_0 ({10'b1011011010, _X_, _X_,
       _X_}), .in_1 ({10'b1011011010, _X_, _X_, _X_}), .in_2
       (13'b0000000110100), .in_3 (13'b1000011100100), .in_4
       (13'b0100000011100), .in_5 (13'b0111000010100), .in_6
       (13'b0111100011100), .in_7 (13'b0000001010100), .in_8
       (13'b0111100010100), .in_9 (13'b0111000010100), .in_10
       (13'b0111100011100), .in_11 (13'b0011101010011), .z ({n_25451,
       n_25443, n_25435, n_25427, n_25419, n_25411, n_25403, n_25395,
       n_25387, n_25379, n_24391, n_24382, n_24373}));
  fx68k_case_box_155 ctl_1310_19(.in_0 (col), .out_0 ({n_24316,
       n_24317, n_24318, n_24319, n_24320, n_24321, n_24322, n_24323,
       n_24324, n_24325, n_24326, n_24327, UNCONNECTED148}));
  fx68k_mux_547 \mux_cmbsop_arA1[3]_1310_19 (.ctl ({n_24316, n_24317,
       n_24318, n_24319, n_24320, n_24321, n_24322, n_24323, n_24324,
       n_24325, n_24326, n_24327}), .in_0 ({10'b0111101011, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_1 ({10'b0111101011, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_2 (17'b00000001101000100), .in_3
       (17'b10000111001000100), .in_4 (17'b01000000111000100), .in_5
       (17'b01110000101000100), .in_6 (17'b01111000111000100), .in_7
       (17'b00000010101000100), .in_8 (17'b01111000101000100), .in_9
       (17'b01110000101000100), .in_10 (17'b01111000111000100), .in_11
       (17'b00111010100111011), .z ({n_25452, n_25444, n_25436,
       n_25428, n_25420, n_25412, n_25404, n_25396, n_25388, n_25380,
       n_24395, n_24392, n_24383, n_24378, n_24374, n_24369, n_24365}));
  fx68k_case_box_158 ctl_1327_19(.in_0 (col), .out_0 ({n_24328,
       n_24329, n_24330, n_24331, n_24332, n_24333, n_24334, n_24335,
       n_24336, n_24337, n_24338, n_24339, UNCONNECTED149}));
  fx68k_mux_520 \mux_cmbsop_arA1[3]_1327_19 (.ctl ({n_24328, n_24329,
       n_24330, n_24331, n_24332, n_24333, n_24334, n_24335, n_24336,
       n_24337, n_24338, n_24339}), .in_0 ({10'b1011011001, _X_, _X_,
       _X_, _X_}), .in_1 ({10'b1011011001, _X_, _X_, _X_, _X_}), .in_2
       (14'b00000001101000), .in_3 (14'b10000111001000), .in_4
       (14'b01000000111000), .in_5 (14'b01110000101000), .in_6
       (14'b01111000111000), .in_7 (14'b00000010101000), .in_8
       (14'b01111000101000), .in_9 (14'b01110000101000), .in_10
       (14'b01111000111000), .in_11 (14'b00111010100111), .z ({n_25453,
       n_25445, n_25437, n_25429, n_25421, n_25413, n_25405, n_25397,
       n_25389, n_25381, n_24393, n_24384, n_24375, n_24366}));
  fx68k_case_box_161 ctl_1344_19(.in_0 (col), .out_0 ({n_24340,
       n_24341, n_24342, n_24343, n_24344, n_24345, n_24346, n_24347,
       n_24348, n_24349, n_24350, n_24351, UNCONNECTED150}));
  fx68k_mux_520 \mux_cmbsop_arA1[3]_1344_19 (.ctl ({n_24340, n_24341,
       n_24342, n_24343, n_24344, n_24345, n_24346, n_24347, n_24348,
       n_24349, n_24350, n_24351}), .in_0 ({10'b0111101010, _X_, _X_,
       _X_, _X_}), .in_1 ({10'b0111101010, _X_, _X_, _X_, _X_}), .in_2
       (14'b00000001101001), .in_3 (14'b10000111001001), .in_4
       (14'b01000000111001), .in_5 (14'b01110000101001), .in_6
       (14'b01111000111001), .in_7 (14'b00000010101001), .in_8
       (14'b01111000101001), .in_9 (14'b01110000101001), .in_10
       (14'b01111000111001), .in_11 (14'b00111010100110), .z ({n_25454,
       n_25446, n_25438, n_25430, n_25422, n_25414, n_25406, n_25398,
       n_25390, n_25382, n_24396, n_24386, n_24385, n_24367}));
  fx68k_mux_671 \mux_arA23[3]_1205_14 (.ctl ({n_24352, n_24353,
       n_24354, n_24355, n_24356, n_24357, n_24358, n_24359, n_24360}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b1), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .z (\arA23[3] [2]));
  fx68k_bmux_546 \mux_arA23[3]_1205_24 (.ctl (movEa), .in_0
       ({\cmbsop_arA1[3] [9], \cmbsop_arA1[3] [8], \cmbsop_arA1[3] [7],
       1'b0, \cmbsop_arA1[3] [5], \cmbsop_arA1[3] [4],
       \cmbsop_arA1[3] [3], \cmbsop_arA1[3] [1], 1'b1}), .in_1
       ({n_24394, n_24387, 2'b01, n_24376, 3'b110, n_24361}), .in_2
       ({1'b1, n_24388, 1'b1, n_24379, 1'b1, n_24370, 2'b11, n_24362}),
       .in_3 ({1'b1, n_24389, 1'b1, n_24380, 1'b1, n_24371, 2'b11,
       n_24363}), .in_4 ({1'b1, n_24390, 1'b1, n_24381, n_24377,
       n_24372, 1'b1, n_24368, n_24364}), .in_5 ({1'b1, n_24391, 1'b1,
       n_24382, 1'b0, n_24373, 3'b110}), .in_6 ({n_24395, n_24392,
       1'b1, n_24383, n_24378, n_24374, 1'b1, n_24369, n_24365}), .in_7
       ({1'b1, n_24393, 1'b1, n_24384, 1'b0, n_24375, 2'b10, n_24366}),
       .in_8 ({n_24396, 1'b1, n_24386, n_24385, 4'b1011, n_24367}), .z
       ({\arA23[3] [9], \arA23[3] [8], \arA23[3] [7], \arA23[3] [6],
       \arA23[3] [5], \arA23[3] [4], \arA23[3] [3], \arA23[3] [1],
       \arA23[3] [0]}));
  fx68k_case_box_167 ctl_548_19(.in_0 (col), .out_0 ({n_24397,
       UNCONNECTED155, n_24398, n_24399, n_24400, n_24401, n_24402,
       n_24403, n_24404, UNCONNECTED154, UNCONNECTED153,
       UNCONNECTED152, UNCONNECTED151}));
  fx68k_mux_93 \mux_cmbsop_arA1[4]_548_19 (.ctl ({n_24397, n_24398,
       n_24399, n_24400, n_24401, n_24402, n_24403, n_24404}), .in_0
       (10'b0100110011), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z
       ({\cmbsop_arA1[4] [19], \cmbsop_arA1[4] [18],
       \cmbsop_arA1[4] [17], \cmbsop_arA1[4] [16], \cmbsop_arA1[4]
       [15], \cmbsop_arA1[4] [14], \cmbsop_arA1[4] [13],
       \cmbsop_arA1[4] [12], \cmbsop_arA1[4] [11], \cmbsop_arA1[4]
       [10]}));
  fx68k_case_box_170 ctl_566_19(.in_0 (col), .out_0 ({n_24405,
       UNCONNECTED160, n_24406, n_24407, n_24408, n_24409, n_24410,
       n_24411, n_24412, UNCONNECTED159, UNCONNECTED158,
       UNCONNECTED157, UNCONNECTED156}));
  fx68k_mux_93 \mux_cmbsop_arA1[4]_566_19 (.ctl ({n_24405, n_24406,
       n_24407, n_24408, n_24409, n_24410, n_24411, n_24412}), .in_0
       (10'b0100110011), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_25732, n_25729,
       n_25726, n_25723, n_25720, n_25717, n_25714, n_25711, n_25708,
       n_25705}));
  fx68k_case_box_173 ctl_584_19(.in_0 (col), .out_0 ({n_24413,
       UNCONNECTED165, n_24414, n_24415, n_24416, n_24417, n_24418,
       n_24419, n_24420, UNCONNECTED164, UNCONNECTED163,
       UNCONNECTED162, UNCONNECTED161}));
  fx68k_mux_77 \mux_cmbsop_arA1[4]_584_19 (.ctl ({n_24413, n_24414,
       n_24415, n_24416, n_24417, n_24418, n_24419, n_24420}), .in_0
       (9'b100110111), .in_1 (9'b000001011), .in_2 (9'b000001111),
       .in_3 (9'b101111001), .in_4 (9'b111000110), .in_5
       (9'b111100111), .in_6 (9'b000001110), .in_7 (9'b111100110), .z
       ({n_25730, n_25727, n_25724, n_25721, n_25718, n_25715, n_25712,
       n_25709, n_25706}));
  fx68k_case_box_176 ctl_602_19(.in_0 (col), .out_0 ({n_24421,
       UNCONNECTED170, n_24422, n_24423, n_24424, n_24425, n_24426,
       n_24427, n_24428, UNCONNECTED169, UNCONNECTED168,
       UNCONNECTED167, UNCONNECTED166}));
  fx68k_mux_93 \mux_cmbsop_arA1[4]_602_19 (.ctl ({n_24421, n_24422,
       n_24423, n_24424, n_24425, n_24426, n_24427, n_24428}), .in_0
       (10'b1110100101), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_25694, n_25684,
       n_25672, n_25661, n_25651, n_25639, n_25627, n_25615, n_25603,
       n_25591}));
  fx68k_case_box_179 ctl_620_19(.in_0 (col), .out_0 ({n_24429,
       UNCONNECTED172, n_24430, n_24431, n_24432, n_24433, n_24434,
       n_24435, n_24436, n_24437, n_24438, n_24439, UNCONNECTED171}));
  fx68k_mux_320 \mux_cmbsop_arA1[4]_620_19 (.ctl ({n_24429, n_24430,
       n_24431, n_24432, n_24433, n_24434, n_24435, n_24436, n_24437,
       n_24438, n_24439}), .in_0 ({10'b1100000001, _X_, _X_, _X_,
       _X_}), .in_1 (14'b00000001100111), .in_2 (14'b10000111000111),
       .in_3 (14'b01000000110111), .in_4 (14'b01110000100111), .in_5
       (14'b01111000110111), .in_6 (14'b00000010100111), .in_7
       (14'b01111000100111), .in_8 (14'b01110000100111), .in_9
       (14'b01111000110111), .in_10 (14'b00111010101000), .z ({n_25695,
       n_25685, n_25673, n_25662, n_25652, n_25640, n_25628, n_25616,
       n_25604, n_25592, n_24528, n_24526, n_24524, n_24522}));
  fx68k_case_box_182 ctl_638_19(.in_0 (col), .out_0 ({n_24440,
       UNCONNECTED174, n_24441, n_24442, n_24443, n_24444, n_24445,
       n_24446, n_24447, n_24448, n_24449, n_24450, UNCONNECTED173}));
  fx68k_mux_320 \mux_cmbsop_arA1[4]_638_19 (.ctl ({n_24440, n_24441,
       n_24442, n_24443, n_24444, n_24445, n_24446, n_24447, n_24448,
       n_24449, n_24450}), .in_0 ({10'b1100000001, _X_, _X_, _X_,
       _X_}), .in_1 (14'b00000001100111), .in_2 (14'b10000111000111),
       .in_3 (14'b01000000110111), .in_4 (14'b01110000100111), .in_5
       (14'b01111000110111), .in_6 (14'b00000010100111), .in_7
       (14'b01111000100111), .in_8 (14'b01110000100111), .in_9
       (14'b01111000110111), .in_10 (14'b00111010101000), .z ({n_25696,
       n_25686, n_25674, n_25663, n_25653, n_25641, n_25629, n_25617,
       n_25605, n_25593, n_24529, n_24527, n_24525, n_24523}));
  fx68k_case_box_185 ctl_656_19(.in_0 (col), .out_0 ({n_24451,
       UNCONNECTED179, n_24452, n_24453, n_24454, n_24455, n_24456,
       n_24457, n_24458, UNCONNECTED178, UNCONNECTED177,
       UNCONNECTED176, UNCONNECTED175}));
  fx68k_mux_93 \mux_cmbsop_arA1[4]_656_19 (.ctl ({n_24451, n_24452,
       n_24453, n_24454, n_24455, n_24456, n_24457, n_24458}), .in_0
       (10'b0100111011), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_25697, n_25687,
       n_25675, n_25664, n_25654, n_25642, n_25630, n_25618, n_25606,
       n_25594}));
  fx68k_case_box_188 ctl_728_19(.in_0 (col), .out_0 ({n_24459,
       UNCONNECTED184, n_24460, n_24461, n_24462, n_24463, n_24464,
       n_24465, n_24466, UNCONNECTED183, UNCONNECTED182,
       UNCONNECTED181, UNCONNECTED180}));
  fx68k_mux_93 \mux_cmbsop_arA1[4]_728_19 (.ctl ({n_24459, n_24460,
       n_24461, n_24462, n_24463, n_24464, n_24465, n_24466}), .in_0
       (10'b0100101101), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_25701, n_25689,
       n_25679, n_25667, n_25656, n_25646, n_25634, n_25622, n_25610,
       n_25598}));
  fx68k_case_box_191 ctl_746_19(.in_0 (col), .out_0 ({n_24467,
       UNCONNECTED189, n_24468, n_24469, n_24470, n_24471, n_24472,
       n_24473, n_24474, UNCONNECTED188, UNCONNECTED187,
       UNCONNECTED186, UNCONNECTED185}));
  fx68k_mux_93 \mux_cmbsop_arA1[4]_746_19 (.ctl ({n_24467, n_24468,
       n_24469, n_24470, n_24471, n_24472, n_24473, n_24474}), .in_0
       (10'b0100101101), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_25702, n_25690,
       n_25680, n_25668, n_25657, n_25647, n_25635, n_25623, n_25611,
       n_25599}));
  fx68k_case_box_194 ctl_764_19(.in_0 (col), .out_0 ({n_24475,
       UNCONNECTED194, n_24476, n_24477, n_24478, n_24479, n_24480,
       n_24481, n_24482, UNCONNECTED193, UNCONNECTED192,
       UNCONNECTED191, UNCONNECTED190}));
  fx68k_mux_77 \mux_cmbsop_arA1[4]_764_19 (.ctl ({n_24475, n_24476,
       n_24477, n_24478, n_24479, n_24480, n_24481, n_24482}), .in_0
       (9'b100100101), .in_1 (9'b000001011), .in_2 (9'b000001111),
       .in_3 (9'b101111001), .in_4 (9'b111000110), .in_5
       (9'b111100111), .in_6 (9'b000001110), .in_7 (9'b111100110), .z
       ({n_25691, n_25681, n_25669, n_25658, n_25648, n_25636, n_25624,
       n_25612, n_25600}));
  fx68k_case_box_197 ctl_782_19(.in_0 (col), .out_0 ({n_24483,
       UNCONNECTED199, n_24484, n_24485, n_24486, n_24487, n_24488,
       n_24489, n_24490, UNCONNECTED198, UNCONNECTED197,
       UNCONNECTED196, UNCONNECTED195}));
  fx68k_mux_93 \mux_cmbsop_arA1[4]_782_19 (.ctl ({n_24483, n_24484,
       n_24485, n_24486, n_24487, n_24488, n_24489, n_24490}), .in_0
       (10'b1101000101), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_25703, n_25692,
       n_25682, n_25670, n_25659, n_25649, n_25637, n_25625, n_25613,
       n_25601}));
  fx68k_case_box_200 ctl_800_19(.in_0 (col), .out_0 ({UNCONNECTED204,
       UNCONNECTED203, n_24492, n_24493, UNCONNECTED202, n_24494,
       n_24495, n_24496, n_24497, n_24498, n_24499, UNCONNECTED201,
       UNCONNECTED200}));
  fx68k_mux_778 \mux_cmbsop_arA1[4]_800_19 (.ctl ({n_24492, n_24493,
       n_24494, n_24495, n_24496, n_24497, n_24498, n_24499}), .in_0
       (16'b0000110000000000), .in_1 (16'b0000010000000000), .in_2
       (16'b1111100000000000), .in_3 (16'b1110100000000000), .in_4
       (16'b1111000000000000), .in_5 (16'b1101000000000000), .in_6
       (16'b1111100000000000), .in_7 (16'b1110100000000000), .z
       ({n_25584, n_25582, n_25579, n_25577, n_25575, n_25573,
       UNCONNECTED214, UNCONNECTED213, UNCONNECTED212, UNCONNECTED211,
       UNCONNECTED210, UNCONNECTED209, UNCONNECTED208, UNCONNECTED207,
       UNCONNECTED206, UNCONNECTED205}));
  fx68k_case_box_203 ctl_818_19(.in_0 (col), .out_0 ({n_24500,
       UNCONNECTED216, n_24501, n_24502, n_24503, n_24504, n_24505,
       n_24506, n_24507, n_24508, n_24509, n_24510, UNCONNECTED215}));
  fx68k_mux_793 \mux_cmbsop_arA1[4]_818_19 (.ctl ({n_24500, n_24501,
       n_24502, n_24503, n_24504, n_24505, n_24506, n_24507, n_24508,
       n_24509, n_24510}), .in_0 ({10'b0101010010, _X_, _X_}), .in_1
       (12'b000000011001), .in_2 (12'b100001110001), .in_3
       (12'b010000001101), .in_4 (12'b011100001001), .in_5
       (12'b011110001101), .in_6 (12'b000000101001), .in_7
       (12'b011110001001), .in_8 (12'b011100001001), .in_9
       (12'b011110001101), .in_10 (12'b001110101010), .z ({n_25569,
       n_25566, n_25563, n_25561, n_25559, n_25556, n_25553, n_25550,
       n_25547, n_25544, n_24521, n_24520}));
  fx68k_mux_804 \mux_arA23[4]_601_10 (.ctl ({n_24511, n_24512, n_24513,
       n_24514, n_24515, n_24516, n_24517, n_24518, n_24519}), .in_0
       (9'b110100001), .in_1 ({n_24528, 1'b0, n_24526, 1'b0, n_24524,
       n_24522, 3'b001}), .in_2 ({n_24529, 1'b0, n_24527, 1'b0,
       n_24525, n_24523, 3'b001}), .in_3 (9'b001011100), .in_4
       (9'b111000011), .in_5 (9'b111000011), .in_6 (9'b111001011),
       .in_7 (9'b101000011), .in_8 ({7'b0010100, n_24521, n_24520}), .z
       ({n_24548, n_24547, n_24546, n_24545, n_24544, n_24543, n_24542,
       n_24541, n_24540}));
  fx68k_mux_812 \mux_arA23[4]_547_19 (.ctl ({n_24536, n_24537, n_24538,
       n_24539}), .in_0 (10'b1010111000), .in_1 (10'b1010111000), .in_2
       (10'b1010111100), .in_3 ({n_24548, 1'b1, n_24547, n_24546,
       n_24545, n_24544, n_24543, n_24542, n_24541, n_24540}), .z
       ({\arA23[4] [9], \arA23[4] [8], \arA23[4] [7], \arA23[4] [6],
       \arA23[4] [5], \arA23[4] [4], \arA23[4] [3], \arA23[4] [2],
       \arA23[4] [1], \arA23[4] [0]}));
  fx68k_case_box_212 ctl_1368_19(.in_0 (col), .out_0 ({n_24549,
       UNCONNECTED218, n_24550, n_24551, n_24552, n_24553, n_24554,
       n_24555, n_24556, UNCONNECTED217}));
  fx68k_mux_93 \mux_cmbsop_arA1[5]_1368_19 (.ctl ({n_24549, n_24550,
       n_24551, n_24552, n_24553, n_24554, n_24555, n_24556}), .in_0
       (10'b1011011000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z
       ({\cmbsop_arA1[5] [19], \cmbsop_arA1[5] [18],
       \cmbsop_arA1[5] [17], \cmbsop_arA1[5] [16], \cmbsop_arA1[5]
       [15], \cmbsop_arA1[5] [14], \cmbsop_arA1[5] [13],
       \cmbsop_arA1[5] [12], \cmbsop_arA1[5] [11], \cmbsop_arA1[5]
       [10]}));
  fx68k_case_box_215 ctl_1382_19(.in_0 (col), .out_0 ({n_24557,
       n_24558, n_24559, n_24560, n_24561, n_24562, n_24563, n_24564,
       n_24565, UNCONNECTED219}));
  fx68k_mux_41 \mux_cmbsop_arA1[5]_1382_19 (.ctl ({n_24557, n_24558,
       n_24559, n_24560, n_24561, n_24562, n_24563, n_24564, n_24565}),
       .in_0 (10'b1011011000), .in_1 (10'b1011011100), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_25797, n_25790, n_25783, n_25776,
       n_25769, n_25762, n_25755, n_25748, n_25741, n_25734}));
  fx68k_case_box_218 ctl_1396_19(.in_0 (col), .out_0 ({n_24566,
       n_24567, n_24568, n_24569, n_24570, n_24571, n_24572, n_24573,
       n_24574, UNCONNECTED220}));
  fx68k_mux_41 \mux_cmbsop_arA1[5]_1396_19 (.ctl ({n_24566, n_24567,
       n_24568, n_24569, n_24570, n_24571, n_24572, n_24573, n_24574}),
       .in_0 (10'b1011011100), .in_1 (10'b1011011100), .in_2
       (10'b0000001011), .in_3 (10'b0000001111), .in_4
       (10'b0101111001), .in_5 (10'b0111000110), .in_6
       (10'b0111100111), .in_7 (10'b0000001110), .in_8
       (10'b0111100110), .z ({n_25798, n_25791, n_25784, n_25777,
       n_25770, n_25763, n_25756, n_25749, n_25742, n_25735}));
  fx68k_case_box_221 ctl_1410_19(.in_0 (col), .out_0 ({n_24575,
       n_24576, n_24577, n_24578, n_24579, n_24580, n_24581, n_24582,
       n_24583, UNCONNECTED221}));
  fx68k_mux_41 \mux_cmbsop_arA1[5]_1410_19 (.ctl ({n_24575, n_24576,
       n_24577, n_24578, n_24579, n_24580, n_24581, n_24582, n_24583}),
       .in_0 (10'b1110000100), .in_1 (10'b0001101100), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_25799, n_25792, n_25785, n_25778,
       n_25771, n_25764, n_25757, n_25750, n_25743, n_25736}));
  fx68k_case_box_224 ctl_1424_19(.in_0 (col), .out_0 ({n_24584,
       UNCONNECTED223, n_24585, n_24586, n_24587, n_24588, n_24589,
       n_24590, n_24591, UNCONNECTED222}));
  fx68k_mux_93 \mux_cmbsop_arA1[5]_1424_19 (.ctl ({n_24584, n_24585,
       n_24586, n_24587, n_24588, n_24589, n_24590, n_24591}), .in_0
       (10'b1011011000), .in_1 (10'b0000000110), .in_2
       (10'b1000011100), .in_3 (10'b0100000011), .in_4
       (10'b0111000010), .in_5 (10'b0111100011), .in_6
       (10'b0000001010), .in_7 (10'b0111100010), .z ({n_25800, n_25793,
       n_25786, n_25779, n_25772, n_25765, n_25758, n_25751, n_25744,
       n_25737}));
  fx68k_case_box_227 ctl_1438_19(.in_0 (col), .out_0 ({n_24592,
       n_24593, n_24594, n_24595, n_24596, n_24597, n_24598, n_24599,
       n_24600, UNCONNECTED224}));
  fx68k_mux_41 \mux_cmbsop_arA1[5]_1438_19 (.ctl ({n_24592, n_24593,
       n_24594, n_24595, n_24596, n_24597, n_24598, n_24599, n_24600}),
       .in_0 (10'b1011011000), .in_1 (10'b1011011100), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_25801, n_25794, n_25787, n_25780,
       n_25773, n_25766, n_25759, n_25752, n_25745, n_25738}));
  fx68k_case_box_230 ctl_1452_19(.in_0 (col), .out_0 ({n_24601,
       n_24602, n_24603, n_24604, n_24605, n_24606, n_24607, n_24608,
       n_24609, UNCONNECTED225}));
  fx68k_mux_41 \mux_cmbsop_arA1[5]_1452_19 (.ctl ({n_24601, n_24602,
       n_24603, n_24604, n_24605, n_24606, n_24607, n_24608, n_24609}),
       .in_0 (10'b1011011100), .in_1 (10'b1011011100), .in_2
       (10'b0000001011), .in_3 (10'b0000001111), .in_4
       (10'b0101111001), .in_5 (10'b0111000110), .in_6
       (10'b0111100111), .in_7 (10'b0000001110), .in_8
       (10'b0111100110), .z ({n_25802, n_25795, n_25788, n_25781,
       n_25774, n_25767, n_25760, n_25753, n_25746, n_25739}));
  fx68k_case_box_233 ctl_1466_19(.in_0 (col), .out_0 ({n_24610,
       n_24611, n_24612, n_24613, n_24614, n_24615, n_24616, n_24617,
       n_24618, UNCONNECTED226}));
  fx68k_mux_41 \mux_cmbsop_arA1[5]_1466_19 (.ctl ({n_24610, n_24611,
       n_24612, n_24613, n_24614, n_24615, n_24616, n_24617, n_24618}),
       .in_0 (10'b1110000100), .in_1 (10'b0001101100), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_25803, n_25796, n_25789, n_25782,
       n_25775, n_25768, n_25761, n_25754, n_25747, n_25740}));
  fx68k_mux_893 \mux_arA23[5]_1365_14 (.ctl ({n_24619, n_24620,
       n_24621, n_24622, n_41, n_83, n_167, n_125}), .in_0
       (7'b0111011), .in_1 (7'b0111011), .in_2 (7'b0111111), .in_3
       (7'b1000000), .in_4 (7'b0111011), .in_5 (7'b0111011), .in_6
       (7'b0111111), .in_7 (7'b1000000), .z ({\arA23[5] [8],
       \arA23[5] [6], \arA23[5] [5], \arA23[5] [4], \arA23[5] [2],
       \arA23[5] [1], \arA23[5] [0]}));
  fx68k_case_box_239 ctl_1486_19(.in_0 (col), .out_0 ({n_24627,
       UNCONNECTED228, n_24628, n_24629, n_24630, n_24631, n_24632,
       n_24633, n_24634, n_24635, n_24636, n_24637, UNCONNECTED227}));
  fx68k_mux_899 \mux_cmbsop_arA1[8]_1486_19 (.ctl ({n_24627, n_24628,
       n_24629, n_24630, n_24631, n_24632, n_24633, n_24634, n_24635,
       n_24636, n_24637}), .in_0 ({10'b0111000001, _X_}), .in_1
       (11'b00000001101), .in_2 (11'b10000111001), .in_3
       (11'b01000000111), .in_4 (11'b01110000101), .in_5
       (11'b01111000111), .in_6 (11'b00000010101), .in_7
       (11'b01111000101), .in_8 (11'b01110000101), .in_9
       (11'b01111000111), .in_10 (11'b00111010100), .z
       ({\cmbsop_arA1[8] [19], \cmbsop_arA1[8] [18],
       \cmbsop_arA1[8] [17], \cmbsop_arA1[8] [16], \cmbsop_arA1[8]
       [15], \cmbsop_arA1[8] [14], \cmbsop_arA1[8] [13],
       \cmbsop_arA1[8] [12], \cmbsop_arA1[8] [11], \cmbsop_arA1[8]
       [10], \cmbsop_arA1[8] [1]}));
  fx68k_case_box_242 ctl_1503_19(.in_0 (col), .out_0 ({n_24638,
       UNCONNECTED230, n_24639, n_24640, n_24641, n_24642, n_24643,
       n_24644, n_24645, n_24646, n_24647, n_24648, UNCONNECTED229}));
  fx68k_mux_899 \mux_cmbsop_arA1[8]_1503_19 (.ctl ({n_24638, n_24639,
       n_24640, n_24641, n_24642, n_24643, n_24644, n_24645, n_24646,
       n_24647, n_24648}), .in_0 ({10'b0111000001, _X_}), .in_1
       (11'b00000001101), .in_2 (11'b10000111001), .in_3
       (11'b01000000111), .in_4 (11'b01110000101), .in_5
       (11'b01111000111), .in_6 (11'b00000010101), .in_7
       (11'b01111000101), .in_8 (11'b01110000101), .in_9
       (11'b01111000111), .in_10 (11'b00111010100), .z ({n_25875,
       n_25868, n_25861, n_25854, n_25847, n_25840, n_25833, n_25826,
       n_25819, n_25812, n_24713}));
  fx68k_case_box_245 ctl_1520_19(.in_0 (col), .out_0 ({n_24649,
       UNCONNECTED232, n_24650, n_24651, n_24652, n_24653, n_24654,
       n_24655, n_24656, n_24657, n_24658, n_24659, UNCONNECTED231}));
  fx68k_mux_793 \mux_cmbsop_arA1[8]_1520_19 (.ctl ({n_24649, n_24650,
       n_24651, n_24652, n_24653, n_24654, n_24655, n_24656, n_24657,
       n_24658, n_24659}), .in_0 ({9'b111000101, _X_, _X_, _X_}), .in_1
       (12'b000001011101), .in_2 (12'b000001111101), .in_3
       (12'b101111001101), .in_4 (12'b111000110101), .in_5
       (12'b111100111101), .in_6 (12'b000001110101), .in_7
       (12'b111100110101), .in_8 (12'b111000110101), .in_9
       (12'b111100111101), .in_10 (12'b010100111010), .z ({n_25869,
       n_25862, n_25855, n_25848, n_25841, n_25834, n_25827, n_25820,
       n_25813, n_24718, n_24717, n_24714}));
  fx68k_case_box_248 ctl_1537_19(.in_0 (col), .out_0 ({n_24660,
       UNCONNECTED234, n_24661, n_24662, n_24663, n_24664, n_24665,
       n_24666, n_24667, n_24668, n_24669, n_24670, UNCONNECTED233}));
  fx68k_mux_899 \mux_cmbsop_arA1[8]_1537_19 (.ctl ({n_24660, n_24661,
       n_24662, n_24663, n_24664, n_24665, n_24666, n_24667, n_24668,
       n_24669, n_24670}), .in_0 ({10'b0010100110, _X_}), .in_1
       (11'b00000001100), .in_2 (11'b10000111000), .in_3
       (11'b01000000110), .in_4 (11'b01110000100), .in_5
       (11'b01111000110), .in_6 (11'b00000010100), .in_7
       (11'b01111000100), .in_8 (11'b01110000100), .in_9
       (11'b01111000110), .in_10 (11'b00111010101), .z ({n_25876,
       n_25870, n_25863, n_25856, n_25849, n_25842, n_25835, n_25828,
       n_25821, n_25814, n_24715}));
  fx68k_case_box_251 ctl_1554_19(.in_0 (col), .out_0 ({n_24671,
       n_24672, n_24673, n_24674, n_24675, n_24676, n_24677, n_24678,
       n_24679, UNCONNECTED238, UNCONNECTED237, UNCONNECTED236,
       UNCONNECTED235}));
  fx68k_mux_41 \mux_cmbsop_arA1[8]_1554_19 (.ctl ({n_24671, n_24672,
       n_24673, n_24674, n_24675, n_24676, n_24677, n_24678, n_24679}),
       .in_0 (10'b0111001101), .in_1 (10'b0100000111), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_25877, n_25871, n_25864, n_25857,
       n_25850, n_25843, n_25836, n_25829, n_25822, n_25815}));
  fx68k_case_box_254 ctl_1571_19(.in_0 (col), .out_0 ({UNCONNECTED244,
       UNCONNECTED243, n_24680, n_24681, n_24682, n_24683, n_24684,
       n_24685, n_24686, UNCONNECTED242, UNCONNECTED241,
       UNCONNECTED240, UNCONNECTED239}));
  fx68k_mux_272 \mux_cmbsop_arA1[8]_1571_19 (.ctl ({n_24680, n_24681,
       n_24682, n_24683, n_24684, n_24685, n_24686}), .in_0
       (10'b0000000110), .in_1 (10'b1000011100), .in_2
       (10'b0100000011), .in_3 (10'b0111000010), .in_4
       (10'b0111100011), .in_5 (10'b0000001010), .in_6
       (10'b0111100010), .z ({n_25878, n_25872, n_25865, n_25858,
       n_25851, n_25844, n_25837, n_25830, n_25823, n_25816}));
  fx68k_case_box_257 ctl_1588_19(.in_0 (col), .out_0 ({UNCONNECTED250,
       UNCONNECTED249, n_24687, n_24688, n_24689, n_24690, n_24691,
       n_24692, n_24693, UNCONNECTED248, UNCONNECTED247,
       UNCONNECTED246, UNCONNECTED245}));
  fx68k_mux_958 \mux_cmbsop_arA1[8]_1588_19 (.ctl ({n_24687, n_24688,
       n_24689, n_24690, n_24691, n_24692, n_24693}), .in_0
       (9'b000001011), .in_1 (9'b000001111), .in_2 (9'b101111001),
       .in_3 (9'b111000110), .in_4 (9'b111100111), .in_5
       (9'b000001110), .in_6 (9'b111100110), .z ({n_25873, n_25866,
       n_25859, n_25852, n_25845, n_25838, n_25831, n_25824, n_25817}));
  fx68k_case_box_260 ctl_1605_19(.in_0 (col), .out_0 ({n_24694,
       UNCONNECTED252, n_24695, n_24696, n_24697, n_24698, n_24699,
       n_24700, n_24701, n_24702, n_24703, n_24704, UNCONNECTED251}));
  fx68k_mux_899 \mux_cmbsop_arA1[8]_1605_19 (.ctl ({n_24694, n_24695,
       n_24696, n_24697, n_24698, n_24699, n_24700, n_24701, n_24702,
       n_24703, n_24704}), .in_0 ({10'b0010101110, _X_}), .in_1
       (11'b00000001100), .in_2 (11'b10000111000), .in_3
       (11'b01000000110), .in_4 (11'b01110000100), .in_5
       (11'b01111000110), .in_6 (11'b00000010100), .in_7
       (11'b01111000100), .in_8 (11'b01110000100), .in_9
       (11'b01111000110), .in_10 (11'b00111010101), .z ({n_25879,
       n_25874, n_25867, n_25860, n_25853, n_25846, n_25839, n_25832,
       n_25825, n_25818, n_24716}));
  fx68k_mux_976 \mux_arA23[8]_1483_14 (.ctl ({n_24619, n_24620,
       n_24621, n_24622, n_41, n_83, n_167, n_125}), .in_0 (6'b011001),
       .in_1 (6'b011001), .in_2 (6'b011001), .in_3 (6'b000100), .in_4
       (6'b100011), .in_5 (6'b100011), .in_6 (6'b100011), .in_7
       (6'b000100), .z ({\arA23[8] [9], \arA23[8] [8], \arA23[8] [6],
       \arA23[8] [5], \arA23[8] [4], \arA23[8] [0]}));
  fx68k_bmux_981 \mux_arA23[8]_1483_26 (.ctl (opcode[8:6]), .in_0
       ({2'b00, \cmbsop_arA1[8] [1]}), .in_1 ({2'b00, n_24713}), .in_2
       ({n_24718, n_24717, n_24714}), .in_3 ({2'b01, n_24715}), .in_4
       (3'b100), .in_5 (3'b100), .in_6 (3'b110), .in_7 ({2'b11,
       n_24716}), .z ({\arA23[8] [3], \arA23[8] [2], \arA23[8] [1]}));
  fx68k_case_box_266 ctl_1628_19(.in_0 (col), .out_0 ({n_24719,
       UNCONNECTED254, n_24720, n_24721, n_24722, n_24723, n_24724,
       n_24725, n_24726, n_24727, n_24728, n_24729, UNCONNECTED253}));
  fx68k_mux_899 \mux_cmbsop_arA1[9]_1628_19 (.ctl ({n_24719, n_24720,
       n_24721, n_24722, n_24723, n_24724, n_24725, n_24726, n_24727,
       n_24728, n_24729}), .in_0 ({10'b0111000001, _X_}), .in_1
       (11'b00000001101), .in_2 (11'b10000111001), .in_3
       (11'b01000000111), .in_4 (11'b01110000101), .in_5
       (11'b01111000111), .in_6 (11'b00000010101), .in_7
       (11'b01111000101), .in_8 (11'b01110000101), .in_9
       (11'b01111000111), .in_10 (11'b00111010100), .z
       ({\cmbsop_arA1[9] [19], \cmbsop_arA1[9] [18],
       \cmbsop_arA1[9] [17], \cmbsop_arA1[9] [16], \cmbsop_arA1[9]
       [15], \cmbsop_arA1[9] [14], \cmbsop_arA1[9] [13],
       \cmbsop_arA1[9] [12], \cmbsop_arA1[9] [11], \cmbsop_arA1[9]
       [10], \cmbsop_arA1[9] [1]}));
  fx68k_case_box_269 ctl_1645_19(.in_0 (col), .out_0 ({n_24730,
       n_24731, n_24732, n_24733, n_24734, n_24735, n_24736, n_24737,
       n_24738, n_24739, n_24740, n_24741, UNCONNECTED255}));
  fx68k_mux_992 \mux_cmbsop_arA1[9]_1645_19 (.ctl ({n_24730, n_24731,
       n_24732, n_24733, n_24734, n_24735, n_24736, n_24737, n_24738,
       n_24739, n_24740, n_24741}), .in_0 ({10'b0111000001, _X_}),
       .in_1 ({10'b0111000001, _X_}), .in_2 (11'b00000001101), .in_3
       (11'b10000111001), .in_4 (11'b01000000111), .in_5
       (11'b01110000101), .in_6 (11'b01111000111), .in_7
       (11'b00000010101), .in_8 (11'b01111000101), .in_9
       (11'b01110000101), .in_10 (11'b01111000111), .in_11
       (11'b00111010100), .z ({n_25943, n_25936, n_25929, n_25922,
       n_25915, n_25908, n_25901, n_25894, n_25887, n_25880, n_24813}));
  fx68k_case_box_272 ctl_1662_19(.in_0 (col), .out_0 ({n_24742,
       n_24743, n_24744, n_24745, n_24746, n_24747, n_24748, n_24749,
       n_24750, n_24751, n_24752, n_24753, UNCONNECTED256}));
  fx68k_mux_1002 \mux_cmbsop_arA1[9]_1662_19 (.ctl ({n_24742, n_24743,
       n_24744, n_24745, n_24746, n_24747, n_24748, n_24749, n_24750,
       n_24751, n_24752, n_24753}), .in_0 ({9'b111000101, _X_, _X_,
       _X_}), .in_1 ({9'b111000101, _X_, _X_, _X_}), .in_2
       (12'b000001011101), .in_3 (12'b000001111101), .in_4
       (12'b101111001101), .in_5 (12'b111000110101), .in_6
       (12'b111100111101), .in_7 (12'b000001110101), .in_8
       (12'b111100110101), .in_9 (12'b111000110101), .in_10
       (12'b111100111101), .in_11 (12'b010100111010), .z ({n_25937,
       n_25930, n_25923, n_25916, n_25909, n_25902, n_25895, n_25888,
       n_25881, n_24820, n_24817, n_24814}));
  fx68k_case_box_275 ctl_1679_19(.in_0 (col), .out_0 ({n_24754,
       n_24755, n_24756, n_24757, n_24758, n_24759, n_24760, n_24761,
       n_24762, n_24763, n_24764, n_24765, UNCONNECTED257}));
  fx68k_mux_454 \mux_cmbsop_arA1[9]_1679_19 (.ctl ({n_24754, n_24755,
       n_24756, n_24757, n_24758, n_24759, n_24760, n_24761, n_24762,
       n_24763, n_24764, n_24765}), .in_0 ({10'b0111001001, _X_, _X_,
       _X_}), .in_1 ({10'b0111001001, _X_, _X_, _X_}), .in_2
       (13'b0000000110011), .in_3 (13'b1000011100011), .in_4
       (13'b0100000011011), .in_5 (13'b0111000010011), .in_6
       (13'b0111100011011), .in_7 (13'b0000001010011), .in_8
       (13'b0111100010011), .in_9 (13'b0111000010011), .in_10
       (13'b0111100011011), .in_11 (13'b0011101010100), .z ({n_25944,
       n_25938, n_25931, n_25924, n_25917, n_25910, n_25903, n_25896,
       n_25889, n_25882, n_24821, n_24818, n_24815}));
  fx68k_case_box_278 ctl_1696_19(.in_0 (col), .out_0 ({n_24766,
       n_24767, n_24768, n_24769, n_24770, n_24771, n_24772, n_24773,
       n_24774, UNCONNECTED261, UNCONNECTED260, UNCONNECTED259,
       UNCONNECTED258}));
  fx68k_mux_41 \mux_cmbsop_arA1[9]_1696_19 (.ctl ({n_24766, n_24767,
       n_24768, n_24769, n_24770, n_24771, n_24772, n_24773, n_24774}),
       .in_0 (10'b0111000001), .in_1 (10'b0100001111), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_25945, n_25939, n_25932, n_25925,
       n_25918, n_25911, n_25904, n_25897, n_25890, n_25883}));
  fx68k_case_box_281 ctl_1713_19(.in_0 (col), .out_0 ({n_24775,
       n_24776, n_24777, n_24778, n_24779, n_24780, n_24781, n_24782,
       n_24783, UNCONNECTED265, UNCONNECTED264, UNCONNECTED263,
       UNCONNECTED262}));
  fx68k_mux_41 \mux_cmbsop_arA1[9]_1713_19 (.ctl ({n_24775, n_24776,
       n_24777, n_24778, n_24779, n_24780, n_24781, n_24782, n_24783}),
       .in_0 (10'b0111000001), .in_1 (10'b0100001111), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_25946, n_25940, n_25933, n_25926,
       n_25919, n_25912, n_25905, n_25898, n_25891, n_25884}));
  fx68k_case_box_284 ctl_1730_19(.in_0 (col), .out_0 ({n_24784,
       n_24785, n_24786, n_24787, n_24788, n_24789, n_24790, n_24791,
       n_24792, UNCONNECTED269, UNCONNECTED268, UNCONNECTED267,
       UNCONNECTED266}));
  fx68k_mux_804 \mux_cmbsop_arA1[9]_1730_19 (.ctl ({n_24784, n_24785,
       n_24786, n_24787, n_24788, n_24789, n_24790, n_24791, n_24792}),
       .in_0 (9'b111000101), .in_1 (9'b100001011), .in_2
       (9'b000001011), .in_3 (9'b000001111), .in_4 (9'b101111001),
       .in_5 (9'b111000110), .in_6 (9'b111100111), .in_7
       (9'b000001110), .in_8 (9'b111100110), .z ({n_25941, n_25934,
       n_25927, n_25920, n_25913, n_25906, n_25899, n_25892, n_25885}));
  fx68k_case_box_287 ctl_1747_19(.in_0 (col), .out_0 ({n_24793,
       n_24794, n_24795, n_24796, n_24797, n_24798, n_24799, n_24800,
       n_24801, n_24802, n_24803, n_24804, UNCONNECTED270}));
  fx68k_mux_1002 \mux_cmbsop_arA1[9]_1747_19 (.ctl ({n_24793, n_24794,
       n_24795, n_24796, n_24797, n_24798, n_24799, n_24800, n_24801,
       n_24802, n_24803, n_24804}), .in_0 ({9'b111000101, _X_, _X_,
       _X_}), .in_1 ({9'b111000101, _X_, _X_, _X_}), .in_2
       (12'b000001011101), .in_3 (12'b000001111101), .in_4
       (12'b101111001101), .in_5 (12'b111000110101), .in_6
       (12'b111100111101), .in_7 (12'b000001110101), .in_8
       (12'b111100110101), .in_9 (12'b111000110101), .in_10
       (12'b111100111101), .in_11 (12'b010100111010), .z ({n_25942,
       n_25935, n_25928, n_25921, n_25914, n_25907, n_25900, n_25893,
       n_25886, n_24822, n_24819, n_24816}));
  fx68k_mux_1062 \mux_arA23[9]_1625_14 (.ctl ({n_24619, n_24620,
       n_24621, n_24622, n_41, n_83, n_167, n_125}), .in_0 (4'b0110),
       .in_1 (4'b0110), .in_2 (4'b0110), .in_3 (4'b0110), .in_4
       (4'b1001), .in_5 (4'b1001), .in_6 (4'b1001), .in_7 (4'b0110), .z
       ({\arA23[9] [9], \arA23[9] [8], \arA23[9] [6], \arA23[9] [4]}));
  fx68k_bmux_981 \mux_arA23[9]_1625_27 (.ctl (opcode[8:6]), .in_0
       ({2'b00, \cmbsop_arA1[9] [1]}), .in_1 ({2'b00, n_24813}), .in_2
       ({n_24820, n_24817, n_24814}), .in_3 ({n_24821, n_24818,
       n_24815}), .in_4 (3'b100), .in_5 (3'b100), .in_6 (3'b110), .in_7
       ({n_24822, n_24819, n_24816}), .z ({\arA23[9] [3], \arA23[9]
       [2], \arA23[9] [1]}));
  fx68k_case_box_293 ctl_1770_19(.in_0 (col), .out_0 ({n_24823,
       UNCONNECTED272, n_24824, n_24825, n_24826, n_24827, n_24828,
       n_24829, n_24830, n_24831, n_24832, n_24833, UNCONNECTED271}));
  fx68k_mux_899 \mux_cmbsop_arA1[11]_1770_19 (.ctl ({n_24823, n_24824,
       n_24825, n_24826, n_24827, n_24828, n_24829, n_24830, n_24831,
       n_24832, n_24833}), .in_0 ({10'b0111010001, _X_}), .in_1
       (11'b00000001101), .in_2 (11'b10000111001), .in_3
       (11'b01000000111), .in_4 (11'b01110000101), .in_5
       (11'b01111000111), .in_6 (11'b00000010101), .in_7
       (11'b01111000101), .in_8 (11'b01110000101), .in_9
       (11'b01111000111), .in_10 (11'b00111010100), .z
       ({\cmbsop_arA1[11] [19], \cmbsop_arA1[11] [18],
       \cmbsop_arA1[11] [17], \cmbsop_arA1[11] [16],
       \cmbsop_arA1[11] [15], \cmbsop_arA1[11] [14],
       \cmbsop_arA1[11] [13], \cmbsop_arA1[11] [12],
       \cmbsop_arA1[11] [11], \cmbsop_arA1[11] [10],
       \cmbsop_arA1[11] [1]}));
  fx68k_case_box_296 ctl_1787_19(.in_0 (col), .out_0 ({n_24834,
       n_24835, n_24836, n_24837, n_24838, n_24839, n_24840, n_24841,
       n_24842, n_24843, n_24844, n_24845, UNCONNECTED273}));
  fx68k_mux_992 \mux_cmbsop_arA1[11]_1787_19 (.ctl ({n_24834, n_24835,
       n_24836, n_24837, n_24838, n_24839, n_24840, n_24841, n_24842,
       n_24843, n_24844, n_24845}), .in_0 ({10'b0111010001, _X_}),
       .in_1 ({10'b0111010001, _X_}), .in_2 (11'b00000001101), .in_3
       (11'b10000111001), .in_4 (11'b01000000111), .in_5
       (11'b01110000101), .in_6 (11'b01111000111), .in_7
       (11'b00000010101), .in_8 (11'b01111000101), .in_9
       (11'b01110000101), .in_10 (11'b01111000111), .in_11
       (11'b00111010100), .z ({n_26010, n_26003, n_25996, n_25989,
       n_25982, n_25975, n_25968, n_25961, n_25954, n_25947, n_24917}));
  fx68k_case_box_299 ctl_1804_19(.in_0 (col), .out_0 ({n_24846,
       n_24847, n_24848, n_24849, n_24850, n_24851, n_24852, n_24853,
       n_24854, n_24855, n_24856, n_24857, UNCONNECTED274}));
  fx68k_mux_119 \mux_cmbsop_arA1[11]_1804_19 (.ctl ({n_24846, n_24847,
       n_24848, n_24849, n_24850, n_24851, n_24852, n_24853, n_24854,
       n_24855, n_24856, n_24857}), .in_0 ({9'b111010101, _X_}), .in_1
       ({9'b111010101, _X_}), .in_2 (10'b0000010111), .in_3
       (10'b0000011111), .in_4 (10'b1011110011), .in_5
       (10'b1110001101), .in_6 (10'b1111001111), .in_7
       (10'b0000011101), .in_8 (10'b1111001101), .in_9
       (10'b1110001101), .in_10 (10'b1111001111), .in_11
       (10'b0101001110), .z ({n_26004, n_25997, n_25990, n_25983,
       n_25976, n_25969, n_25962, n_25955, n_25948, n_24918}));
  fx68k_case_box_302 ctl_1821_19(.in_0 (col), .out_0 ({n_24858,
       n_24859, n_24860, n_24861, n_24862, n_24863, n_24864, n_24865,
       n_24866, n_24867, n_24868, n_24869, UNCONNECTED275}));
  fx68k_mux_454 \mux_cmbsop_arA1[11]_1821_19 (.ctl ({n_24858, n_24859,
       n_24860, n_24861, n_24862, n_24863, n_24864, n_24865, n_24866,
       n_24867, n_24868, n_24869}), .in_0 ({10'b0111011001, _X_, _X_,
       _X_}), .in_1 ({10'b0111011001, _X_, _X_, _X_}), .in_2
       (13'b0000000110011), .in_3 (13'b1000011100011), .in_4
       (13'b0100000011011), .in_5 (13'b0111000010011), .in_6
       (13'b0111100011011), .in_7 (13'b0000001010011), .in_8
       (13'b0111100010011), .in_9 (13'b0111000010011), .in_10
       (13'b0111100011011), .in_11 (13'b0011101010100), .z ({n_26011,
       n_26005, n_25998, n_25991, n_25984, n_25977, n_25970, n_25963,
       n_25956, n_25949, n_24922, n_24921, n_24919}));
  fx68k_case_box_305 ctl_1838_19(.in_0 (col), .out_0 ({n_24870,
       n_24871, n_24872, n_24873, n_24874, n_24875, n_24876, n_24877,
       n_24878, UNCONNECTED279, UNCONNECTED278, UNCONNECTED277,
       UNCONNECTED276}));
  fx68k_mux_41 \mux_cmbsop_arA1[11]_1838_19 (.ctl ({n_24870, n_24871,
       n_24872, n_24873, n_24874, n_24875, n_24876, n_24877, n_24878}),
       .in_0 (10'b0100000000), .in_1 (10'b0001101011), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_26012, n_26006, n_25999, n_25992,
       n_25985, n_25978, n_25971, n_25964, n_25957, n_25950}));
  fx68k_case_box_308 ctl_1855_19(.in_0 (col), .out_0 ({n_24879,
       n_24880, n_24881, n_24882, n_24883, n_24884, n_24885, n_24886,
       n_24887, UNCONNECTED283, UNCONNECTED282, UNCONNECTED281,
       UNCONNECTED280}));
  fx68k_mux_41 \mux_cmbsop_arA1[11]_1855_19 (.ctl ({n_24879, n_24880,
       n_24881, n_24882, n_24883, n_24884, n_24885, n_24886, n_24887}),
       .in_0 (10'b0100000000), .in_1 (10'b0001101011), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_26013, n_26007, n_26000, n_25993,
       n_25986, n_25979, n_25972, n_25965, n_25958, n_25951}));
  fx68k_case_box_311 ctl_1872_19(.in_0 (col), .out_0 ({n_24888,
       n_24889, n_24890, n_24891, n_24892, n_24893, n_24894, n_24895,
       n_24896, UNCONNECTED287, UNCONNECTED286, UNCONNECTED285,
       UNCONNECTED284}));
  fx68k_mux_804 \mux_cmbsop_arA1[11]_1872_19 (.ctl ({n_24888, n_24889,
       n_24890, n_24891, n_24892, n_24893, n_24894, n_24895, n_24896}),
       .in_0 (9'b100001100), .in_1 (9'b001101111), .in_2
       (9'b000001011), .in_3 (9'b000001111), .in_4 (9'b101111001),
       .in_5 (9'b111000110), .in_6 (9'b111100111), .in_7
       (9'b000001110), .in_8 (9'b111100110), .z ({n_26008, n_26001,
       n_25994, n_25987, n_25980, n_25973, n_25966, n_25959, n_25952}));
  fx68k_case_box_314 ctl_1889_19(.in_0 (col), .out_0 ({n_24897,
       n_24898, n_24899, n_24900, n_24901, n_24902, n_24903, n_24904,
       n_24905, n_24906, n_24907, n_24908, UNCONNECTED288}));
  fx68k_mux_119 \mux_cmbsop_arA1[11]_1889_19 (.ctl ({n_24897, n_24898,
       n_24899, n_24900, n_24901, n_24902, n_24903, n_24904, n_24905,
       n_24906, n_24907, n_24908}), .in_0 ({9'b111010101, _X_}), .in_1
       ({9'b111010101, _X_}), .in_2 (10'b0000010111), .in_3
       (10'b0000011111), .in_4 (10'b1011110011), .in_5
       (10'b1110001101), .in_6 (10'b1111001111), .in_7
       (10'b0000011101), .in_8 (10'b1111001101), .in_9
       (10'b1110001101), .in_10 (10'b1111001111), .in_11
       (10'b0101001110), .z ({n_26009, n_26002, n_25995, n_25988,
       n_25981, n_25974, n_25967, n_25960, n_25953, n_24920}));
  fx68k_mux_1062 \mux_arA23[11]_1767_14 (.ctl ({n_24619, n_24620,
       n_24621, n_24622, n_41, n_83, n_167, n_125}), .in_0 (4'b0110),
       .in_1 (4'b0110), .in_2 (4'b0110), .in_3 (4'b0111), .in_4
       (4'b1001), .in_5 (4'b1001), .in_6 (4'b1001), .in_7 (4'b0110), .z
       ({\arA23[11] [9], \arA23[11] [8], \arA23[11] [6], \arA23[11]
       [3]}));
  fx68k_bmux_981 \mux_arA23[11]_1767_28 (.ctl (opcode[8:6]), .in_0
       ({2'b10, \cmbsop_arA1[11] [1]}), .in_1 ({2'b10, n_24917}), .in_2
       ({2'b11, n_24918}), .in_3 ({n_24922, n_24921, n_24919}), .in_4
       (3'b100), .in_5 (3'b100), .in_6 (3'b110), .in_7 ({2'b11,
       n_24920}), .z ({\arA23[11] [4], \arA23[11] [2], \arA23[11]
       [1]}));
  fx68k_case_box_320 ctl_1912_19(.in_0 (col), .out_0 ({n_24923,
       UNCONNECTED290, n_24924, n_24925, n_24926, n_24927, n_24928,
       n_24929, n_24930, n_24931, n_24932, n_24933, UNCONNECTED289}));
  fx68k_mux_899 \mux_cmbsop_arA1[12]_1912_19 (.ctl ({n_24923, n_24924,
       n_24925, n_24926, n_24927, n_24928, n_24929, n_24930, n_24931,
       n_24932, n_24933}), .in_0 ({10'b0111000001, _X_}), .in_1
       (11'b00000001101), .in_2 (11'b10000111001), .in_3
       (11'b01000000111), .in_4 (11'b01110000101), .in_5
       (11'b01111000111), .in_6 (11'b00000010101), .in_7
       (11'b01111000101), .in_8 (11'b01110000101), .in_9
       (11'b01111000111), .in_10 (11'b00111010100), .z
       ({\cmbsop_arA1[12] [19], \cmbsop_arA1[12] [18],
       \cmbsop_arA1[12] [17], \cmbsop_arA1[12] [16],
       \cmbsop_arA1[12] [15], \cmbsop_arA1[12] [14],
       \cmbsop_arA1[12] [13], \cmbsop_arA1[12] [12],
       \cmbsop_arA1[12] [11], \cmbsop_arA1[12] [10],
       \cmbsop_arA1[12] [1]}));
  fx68k_case_box_323 ctl_1929_19(.in_0 (col), .out_0 ({n_24934,
       UNCONNECTED292, n_24935, n_24936, n_24937, n_24938, n_24939,
       n_24940, n_24941, n_24942, n_24943, n_24944, UNCONNECTED291}));
  fx68k_mux_899 \mux_cmbsop_arA1[12]_1929_19 (.ctl ({n_24934, n_24935,
       n_24936, n_24937, n_24938, n_24939, n_24940, n_24941, n_24942,
       n_24943, n_24944}), .in_0 ({10'b0111000001, _X_}), .in_1
       (11'b00000001101), .in_2 (11'b10000111001), .in_3
       (11'b01000000111), .in_4 (11'b01110000101), .in_5
       (11'b01111000111), .in_6 (11'b00000010101), .in_7
       (11'b01111000101), .in_8 (11'b01110000101), .in_9
       (11'b01111000111), .in_10 (11'b00111010100), .z ({n_26077,
       n_26070, n_26063, n_26056, n_26049, n_26042, n_26035, n_26028,
       n_26021, n_26014, n_25014}));
  fx68k_case_box_326 ctl_1946_19(.in_0 (col), .out_0 ({n_24945,
       UNCONNECTED294, n_24946, n_24947, n_24948, n_24949, n_24950,
       n_24951, n_24952, n_24953, n_24954, n_24955, UNCONNECTED293}));
  fx68k_mux_793 \mux_cmbsop_arA1[12]_1946_19 (.ctl ({n_24945, n_24946,
       n_24947, n_24948, n_24949, n_24950, n_24951, n_24952, n_24953,
       n_24954, n_24955}), .in_0 ({9'b111000101, _X_, _X_, _X_}), .in_1
       (12'b000001011101), .in_2 (12'b000001111101), .in_3
       (12'b101111001101), .in_4 (12'b111000110101), .in_5
       (12'b111100111101), .in_6 (12'b000001110101), .in_7
       (12'b111100110101), .in_8 (12'b111000110101), .in_9
       (12'b111100111101), .in_10 (12'b010100111010), .z ({n_26071,
       n_26064, n_26057, n_26050, n_26043, n_26036, n_26029, n_26022,
       n_26015, n_25017, n_25016, n_25015}));
  fx68k_case_box_329 ctl_1963_19(.in_0 (col), .out_0 ({n_24956,
       UNCONNECTED296, n_24957, n_24958, n_24959, n_24960, n_24961,
       n_24962, n_24963, n_24964, n_24965, n_24966, UNCONNECTED295}));
  fx68k_mux_899 \mux_cmbsop_arA1[12]_1963_19 (.ctl ({n_24956, n_24957,
       n_24958, n_24959, n_24960, n_24961, n_24962, n_24963, n_24964,
       n_24965, n_24966}), .in_0 ({10'b0101011011, _X_}), .in_1
       (11'b00000001100), .in_2 (11'b10000111000), .in_3
       (11'b01000000110), .in_4 (11'b01110000100), .in_5
       (11'b01111000110), .in_6 (11'b00000010100), .in_7
       (11'b01111000100), .in_8 (11'b01110000100), .in_9
       (11'b01111000110), .in_10 (11'b00111010101), .z ({n_26078,
       n_26072, n_26065, n_26058, n_26051, n_26044, n_26037, n_26030,
       n_26023, n_26016, n_25012}));
  fx68k_case_box_332 ctl_1980_19(.in_0 (col), .out_0 ({n_24967,
       n_24968, n_24969, n_24970, n_24971, n_24972, n_24973, n_24974,
       n_24975, UNCONNECTED300, UNCONNECTED299, UNCONNECTED298,
       UNCONNECTED297}));
  fx68k_mux_41 \mux_cmbsop_arA1[12]_1980_19 (.ctl ({n_24967, n_24968,
       n_24969, n_24970, n_24971, n_24972, n_24973, n_24974, n_24975}),
       .in_0 (10'b0111001101), .in_1 (10'b0100000111), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_26079, n_26073, n_26066, n_26059,
       n_26052, n_26045, n_26038, n_26031, n_26024, n_26017}));
  fx68k_case_box_335 ctl_1997_19(.in_0 (col), .out_0 ({n_24976,
       n_24977, n_24978, n_24979, n_24980, n_24981, n_24982, n_24983,
       n_24984, UNCONNECTED304, UNCONNECTED303, UNCONNECTED302,
       UNCONNECTED301}));
  fx68k_mux_41 \mux_cmbsop_arA1[12]_1997_19 (.ctl ({n_24976, n_24977,
       n_24978, n_24979, n_24980, n_24981, n_24982, n_24983, n_24984}),
       .in_0 (10'b1111100011), .in_1 (10'b1111100011), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_26080, n_26074, n_26067, n_26060,
       n_26053, n_26046, n_26039, n_26032, n_26025, n_26018}));
  fx68k_case_box_338 ctl_2014_19(.in_0 (col), .out_0 ({UNCONNECTED309,
       n_24985, n_24986, n_24987, n_24988, n_24989, n_24990, n_24991,
       n_24992, UNCONNECTED308, UNCONNECTED307, UNCONNECTED306,
       UNCONNECTED305}));
  fx68k_mux_93 \mux_cmbsop_arA1[12]_2014_19 (.ctl ({n_24985, n_24986,
       n_24987, n_24988, n_24989, n_24990, n_24991, n_24992}), .in_0
       (10'b1111100011), .in_1 (10'b0000001011), .in_2
       (10'b0000001111), .in_3 (10'b0101111001), .in_4
       (10'b0111000110), .in_5 (10'b0111100111), .in_6
       (10'b0000001110), .in_7 (10'b0111100110), .z ({n_26081, n_26075,
       n_26068, n_26061, n_26054, n_26047, n_26040, n_26033, n_26026,
       n_26019}));
  fx68k_case_box_341 ctl_2031_19(.in_0 (col), .out_0 ({n_24993,
       UNCONNECTED311, n_24994, n_24995, n_24996, n_24997, n_24998,
       n_24999, n_25000, n_25001, n_25002, n_25003, UNCONNECTED310}));
  fx68k_mux_899 \mux_cmbsop_arA1[12]_2031_19 (.ctl ({n_24993, n_24994,
       n_24995, n_24996, n_24997, n_24998, n_24999, n_25000, n_25001,
       n_25002, n_25003}), .in_0 ({10'b0101011011, _X_}), .in_1
       (11'b00000001100), .in_2 (11'b10000111000), .in_3
       (11'b01000000110), .in_4 (11'b01110000100), .in_5
       (11'b01111000110), .in_6 (11'b00000010100), .in_7
       (11'b01111000100), .in_8 (11'b01110000100), .in_9
       (11'b01111000110), .in_10 (11'b00111010101), .z ({n_26082,
       n_26076, n_26069, n_26062, n_26055, n_26048, n_26041, n_26034,
       n_26027, n_26020, n_25013}));
  fx68k_mux_1224 \mux_arA23[12]_1909_14 (.ctl ({n_24619, n_24620,
       n_24621, n_24622, n_41, n_83, n_167, n_125}), .in_0 (5'b01110),
       .in_1 (5'b01110), .in_2 (5'b01110), .in_3 (5'b01011), .in_4
       (5'b10101), .in_5 (5'b10101), .in_6 (5'b10101), .in_7
       (5'b01011), .z ({\arA23[12] [9], \arA23[12] [8], \arA23[12] [7],
       \arA23[12] [6], \arA23[12] [4]}));
  fx68k_bmux_1228 \mux_arA23[12]_1909_29 (.ctl (opcode[8:6]), .in_0
       ({2'b00, \cmbsop_arA1[12] [1], 1'b1}), .in_1 ({2'b00, n_25014,
       1'b1}), .in_2 ({n_25017, n_25016, n_25015, 1'b1}), .in_3
       ({3'b101, n_25012}), .in_4 (4'b1001), .in_5 (4'b1001), .in_6
       (4'b1101), .in_7 ({3'b101, n_25013}), .z ({\arA23[12] [3],
       \arA23[12] [2], \arA23[12] [1], \arA23[12] [0]}));
  fx68k_case_box_347 ctl_2054_19(.in_0 (col), .out_0 ({n_25018,
       UNCONNECTED313, n_25019, n_25020, n_25021, n_25022, n_25023,
       n_25024, n_25025, n_25026, n_25027, n_25028, UNCONNECTED312}));
  fx68k_mux_899 \mux_cmbsop_arA1[13]_2054_19 (.ctl ({n_25018, n_25019,
       n_25020, n_25021, n_25022, n_25023, n_25024, n_25025, n_25026,
       n_25027, n_25028}), .in_0 ({10'b0111000001, _X_}), .in_1
       (11'b00000001101), .in_2 (11'b10000111001), .in_3
       (11'b01000000111), .in_4 (11'b01110000101), .in_5
       (11'b01111000111), .in_6 (11'b00000010101), .in_7
       (11'b01111000101), .in_8 (11'b01110000101), .in_9
       (11'b01111000111), .in_10 (11'b00111010100), .z
       ({\cmbsop_arA1[13] [19], \cmbsop_arA1[13] [18],
       \cmbsop_arA1[13] [17], \cmbsop_arA1[13] [16],
       \cmbsop_arA1[13] [15], \cmbsop_arA1[13] [14],
       \cmbsop_arA1[13] [13], \cmbsop_arA1[13] [12],
       \cmbsop_arA1[13] [11], \cmbsop_arA1[13] [10],
       \cmbsop_arA1[13] [1]}));
  fx68k_case_box_350 ctl_2071_19(.in_0 (col), .out_0 ({n_25029,
       n_25030, n_25031, n_25032, n_25033, n_25034, n_25035, n_25036,
       n_25037, n_25038, n_25039, n_25040, UNCONNECTED314}));
  fx68k_mux_992 \mux_cmbsop_arA1[13]_2071_19 (.ctl ({n_25029, n_25030,
       n_25031, n_25032, n_25033, n_25034, n_25035, n_25036, n_25037,
       n_25038, n_25039, n_25040}), .in_0 ({10'b0111000001, _X_}),
       .in_1 ({10'b0111000001, _X_}), .in_2 (11'b00000001101), .in_3
       (11'b10000111001), .in_4 (11'b01000000111), .in_5
       (11'b01110000101), .in_6 (11'b01111000111), .in_7
       (11'b00000010101), .in_8 (11'b01111000101), .in_9
       (11'b01110000101), .in_10 (11'b01111000111), .in_11
       (11'b00111010100), .z ({n_26146, n_26139, n_26132, n_26125,
       n_26118, n_26111, n_26104, n_26097, n_26090, n_26083, n_25112}));
  fx68k_case_box_353 ctl_2088_19(.in_0 (col), .out_0 ({n_25041,
       n_25042, n_25043, n_25044, n_25045, n_25046, n_25047, n_25048,
       n_25049, n_25050, n_25051, n_25052, UNCONNECTED315}));
  fx68k_mux_1002 \mux_cmbsop_arA1[13]_2088_19 (.ctl ({n_25041, n_25042,
       n_25043, n_25044, n_25045, n_25046, n_25047, n_25048, n_25049,
       n_25050, n_25051, n_25052}), .in_0 ({9'b111000101, _X_, _X_,
       _X_}), .in_1 ({9'b111000101, _X_, _X_, _X_}), .in_2
       (12'b000001011101), .in_3 (12'b000001111101), .in_4
       (12'b101111001101), .in_5 (12'b111000110101), .in_6
       (12'b111100111101), .in_7 (12'b000001110101), .in_8
       (12'b111100110101), .in_9 (12'b111000110101), .in_10
       (12'b111100111101), .in_11 (12'b010100111010), .z ({n_26140,
       n_26133, n_26126, n_26119, n_26112, n_26105, n_26098, n_26091,
       n_26084, n_25119, n_25116, n_25113}));
  fx68k_case_box_356 ctl_2105_19(.in_0 (col), .out_0 ({n_25053,
       n_25054, n_25055, n_25056, n_25057, n_25058, n_25059, n_25060,
       n_25061, n_25062, n_25063, n_25064, UNCONNECTED316}));
  fx68k_mux_454 \mux_cmbsop_arA1[13]_2105_19 (.ctl ({n_25053, n_25054,
       n_25055, n_25056, n_25057, n_25058, n_25059, n_25060, n_25061,
       n_25062, n_25063, n_25064}), .in_0 ({10'b0111001001, _X_, _X_,
       _X_}), .in_1 ({10'b0111001001, _X_, _X_, _X_}), .in_2
       (13'b0000000110011), .in_3 (13'b1000011100011), .in_4
       (13'b0100000011011), .in_5 (13'b0111000010011), .in_6
       (13'b0111100011011), .in_7 (13'b0000001010011), .in_8
       (13'b0111100010011), .in_9 (13'b0111000010011), .in_10
       (13'b0111100011011), .in_11 (13'b0011101010100), .z ({n_26147,
       n_26141, n_26134, n_26127, n_26120, n_26113, n_26106, n_26099,
       n_26092, n_26085, n_25120, n_25117, n_25114}));
  fx68k_case_box_359 ctl_2122_19(.in_0 (col), .out_0 ({n_25065,
       n_25066, n_25067, n_25068, n_25069, n_25070, n_25071, n_25072,
       n_25073, UNCONNECTED320, UNCONNECTED319, UNCONNECTED318,
       UNCONNECTED317}));
  fx68k_mux_41 \mux_cmbsop_arA1[13]_2122_19 (.ctl ({n_25065, n_25066,
       n_25067, n_25068, n_25069, n_25070, n_25071, n_25072, n_25073}),
       .in_0 (10'b0111000001), .in_1 (10'b0100001111), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_26148, n_26142, n_26135, n_26128,
       n_26121, n_26114, n_26107, n_26100, n_26093, n_26086}));
  fx68k_case_box_362 ctl_2139_19(.in_0 (col), .out_0 ({n_25074,
       n_25075, n_25076, n_25077, n_25078, n_25079, n_25080, n_25081,
       n_25082, UNCONNECTED324, UNCONNECTED323, UNCONNECTED322,
       UNCONNECTED321}));
  fx68k_mux_41 \mux_cmbsop_arA1[13]_2139_19 (.ctl ({n_25074, n_25075,
       n_25076, n_25077, n_25078, n_25079, n_25080, n_25081, n_25082}),
       .in_0 (10'b0111000001), .in_1 (10'b0100001111), .in_2
       (10'b0000000110), .in_3 (10'b1000011100), .in_4
       (10'b0100000011), .in_5 (10'b0111000010), .in_6
       (10'b0111100011), .in_7 (10'b0000001010), .in_8
       (10'b0111100010), .z ({n_26149, n_26143, n_26136, n_26129,
       n_26122, n_26115, n_26108, n_26101, n_26094, n_26087}));
  fx68k_case_box_365 ctl_2156_19(.in_0 (col), .out_0 ({n_25083,
       n_25084, n_25085, n_25086, n_25087, n_25088, n_25089, n_25090,
       n_25091, UNCONNECTED328, UNCONNECTED327, UNCONNECTED326,
       UNCONNECTED325}));
  fx68k_mux_804 \mux_cmbsop_arA1[13]_2156_19 (.ctl ({n_25083, n_25084,
       n_25085, n_25086, n_25087, n_25088, n_25089, n_25090, n_25091}),
       .in_0 (9'b111000101), .in_1 (9'b100001011), .in_2
       (9'b000001011), .in_3 (9'b000001111), .in_4 (9'b101111001),
       .in_5 (9'b111000110), .in_6 (9'b111100111), .in_7
       (9'b000001110), .in_8 (9'b111100110), .z ({n_26144, n_26137,
       n_26130, n_26123, n_26116, n_26109, n_26102, n_26095, n_26088}));
  fx68k_case_box_368 ctl_2173_19(.in_0 (col), .out_0 ({n_25092,
       n_25093, n_25094, n_25095, n_25096, n_25097, n_25098, n_25099,
       n_25100, n_25101, n_25102, n_25103, UNCONNECTED329}));
  fx68k_mux_1002 \mux_cmbsop_arA1[13]_2173_19 (.ctl ({n_25092, n_25093,
       n_25094, n_25095, n_25096, n_25097, n_25098, n_25099, n_25100,
       n_25101, n_25102, n_25103}), .in_0 ({9'b111000101, _X_, _X_,
       _X_}), .in_1 ({9'b111000101, _X_, _X_, _X_}), .in_2
       (12'b000001011101), .in_3 (12'b000001111101), .in_4
       (12'b101111001101), .in_5 (12'b111000110101), .in_6
       (12'b111100111101), .in_7 (12'b000001110101), .in_8
       (12'b111100110101), .in_9 (12'b111000110101), .in_10
       (12'b111100111101), .in_11 (12'b010100111010), .z ({n_26145,
       n_26138, n_26131, n_26124, n_26117, n_26110, n_26103, n_26096,
       n_26089, n_25121, n_25118, n_25115}));
  fx68k_mux_1062 \mux_arA23[13]_2051_14 (.ctl ({n_24619, n_24620,
       n_24621, n_24622, n_41, n_83, n_167, n_125}), .in_0 (4'b0110),
       .in_1 (4'b0110), .in_2 (4'b0110), .in_3 (4'b0110), .in_4
       (4'b1001), .in_5 (4'b1001), .in_6 (4'b1001), .in_7 (4'b0110), .z
       ({\arA23[13] [9], \arA23[13] [8], \arA23[13] [6], \arA23[13]
       [4]}));
  fx68k_bmux_981 \mux_arA23[13]_2051_30 (.ctl (opcode[8:6]), .in_0
       ({2'b00, \cmbsop_arA1[13] [1]}), .in_1 ({2'b00, n_25112}), .in_2
       ({n_25119, n_25116, n_25113}), .in_3 ({n_25120, n_25117,
       n_25114}), .in_4 (3'b100), .in_5 (3'b100), .in_6 (3'b110), .in_7
       ({n_25121, n_25118, n_25115}), .z ({\arA23[13] [3],
       \arA23[13] [2], \arA23[13] [1]}));
  fx68k_bmux_1313 \mux_arA23[line]_79_40 (.ctl (opcode[15:12]), .in_0
       ({\arA23[0] [9], \arA23[0] [8], \arA23[0] [7], \arA23[0] [6],
       \arA23[0] [5], \arA23[0] [4], \arA23[0] [3], \arA23[0] [2],
       \arA23[0] [1], \arA23[0] [0]}), .in_1 ({\arA23[1] [9],
       \arA23[1] [8], \arA23[1] [7], \arA23[1] [6], \arA23[1] [5],
       \arA23[1] [4], \arA23[1] [3], \arA23[1] [2], \arA23[1] [1],
       \arA23[1] [0]}), .in_2 ({\arA23[2] [9], \arA23[2] [8],
       \arA23[2] [7], \arA23[2] [6], \arA23[2] [5], \arA23[2] [4],
       1'b1, \arA23[2] [2], \arA23[2] [1], \arA23[2] [0]}), .in_3
       ({\arA23[3] [9], \arA23[3] [8], \arA23[3] [7], \arA23[3] [6],
       \arA23[3] [5], \arA23[3] [4], \arA23[3] [3], \arA23[3] [2],
       \arA23[3] [1], \arA23[3] [0]}), .in_4 ({\arA23[4] [9],
       \arA23[4] [8], \arA23[4] [7], \arA23[4] [6], \arA23[4] [5],
       \arA23[4] [4], \arA23[4] [3], \arA23[4] [2], \arA23[4] [1],
       \arA23[4] [0]}), .in_5 ({1'b1, \arA23[5] [8], 1'b1, \arA23[5]
       [6], \arA23[5] [5], \arA23[5] [4], 1'b0, \arA23[5] [2],
       \arA23[5] [1], \arA23[5] [0]}), .in_6 ({_X_, _X_, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_7 ({_X_, _X_, _X_, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_8 ({\arA23[8] [9], \arA23[8] [8],
       1'b1, \arA23[8] [6], \arA23[8] [5], \arA23[8] [4], \arA23[8]
       [3], \arA23[8] [2], \arA23[8] [1], \arA23[8] [0]}), .in_9
       ({\arA23[9] [9], \arA23[9] [8], 1'b1, \arA23[9] [6], 1'b0,
       \arA23[9] [4], \arA23[9] [3], \arA23[9] [2], \arA23[9] [1],
       1'b1}), .in_10 ({_X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_,
       _X_}), .in_11 ({\arA23[11] [9], \arA23[11] [8], 1'b1,
       \arA23[11] [6], 1'b0, \arA23[11] [4], \arA23[11] [3],
       \arA23[11] [2], \arA23[11] [1], 1'b1}), .in_12 ({\arA23[12] [9],
       \arA23[12] [8], \arA23[12] [7], \arA23[12] [6], 1'b0,
       \arA23[12] [4], \arA23[12] [3], \arA23[12] [2], \arA23[12] [1],
       \arA23[12] [0]}), .in_13 ({\arA23[13] [9], \arA23[13] [8], 1'b1,
       \arA23[13] [6], 1'b0, \arA23[13] [4], \arA23[13] [3],
       \arA23[13] [2], \arA23[13] [1], 1'b1}), .in_14 (10'b1111000111),
       .in_15 ({_X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_}), .z
       ({\arA23[line] [9], \arA23[line] [8], \arA23[line] [7],
       \arA23[line] [6], \arA23[line] [5], \arA23[line] [4],
       \arA23[line] [3], \arA23[line] [2], \arA23[line] [1],
       \arA23[line] [0]}));
  fx68k_bmux_299 mux_79_19(.ctl (lineBmap[0]), .in_0 ({\arA23[line]
       [9], \arA23[line] [8], \arA23[line] [7], \arA23[line] [6],
       \arA23[line] [5], \arA23[line] [4], \arA23[line] [3],
       \arA23[line] [2], \arA23[line] [1], \arA23[line] [0]}), .in_1
       ({scA3[9], 1'b0, scA3[7:1], 1'b1}), .z (plaA3));
  fx68k_bmux_1313 \mux_arA23[line]_78_19 (.ctl (opcode[15:12]), .in_0
       ({\arA23[0] [9], \arA23[0] [8], \arA23[0] [7], \arA23[0] [6],
       \arA23[0] [5], \arA23[0] [4], \arA23[0] [3], \arA23[0] [2],
       \arA23[0] [1], \arA23[0] [0]}), .in_1 ({\arA23[1] [9],
       \arA23[1] [8], \arA23[1] [7], \arA23[1] [6], \arA23[1] [5],
       \arA23[1] [4], \arA23[1] [3], \arA23[1] [2], \arA23[1] [1],
       \arA23[1] [0]}), .in_2 ({\arA23[2] [9], \arA23[2] [8],
       \arA23[2] [7], \arA23[2] [6], \arA23[2] [5], \arA23[2] [4],
       1'b1, \arA23[2] [2], \arA23[2] [1], \arA23[2] [0]}), .in_3
       ({\arA23[3] [9], \arA23[3] [8], \arA23[3] [7], \arA23[3] [6],
       \arA23[3] [5], \arA23[3] [4], \arA23[3] [3], \arA23[3] [2],
       \arA23[3] [1], \arA23[3] [0]}), .in_4 ({\arA23[4] [9],
       \arA23[4] [8], \arA23[4] [7], \arA23[4] [6], \arA23[4] [5],
       \arA23[4] [4], \arA23[4] [3], \arA23[4] [2], \arA23[4] [1],
       \arA23[4] [0]}), .in_5 ({1'b1, \arA23[5] [8], 1'b1, \arA23[5]
       [6], \arA23[5] [5], \arA23[5] [4], 1'b0, \arA23[5] [2],
       \arA23[5] [1], \arA23[5] [0]}), .in_6 ({_X_, _X_, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_}), .in_7 ({_X_, _X_, _X_, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_8 ({\arA23[8] [9], \arA23[8] [8],
       1'b1, \arA23[8] [6], \arA23[8] [5], \arA23[8] [4], \arA23[8]
       [3], \arA23[8] [2], \arA23[8] [1], \arA23[8] [0]}), .in_9
       ({\arA23[9] [9], \arA23[9] [8], 1'b1, \arA23[9] [6], 1'b0,
       \arA23[9] [4], \arA23[9] [3], \arA23[9] [2], \arA23[9] [1],
       1'b1}), .in_10 ({_X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_,
       _X_}), .in_11 ({\arA23[11] [9], \arA23[11] [8], 1'b1,
       \arA23[11] [6], 1'b0, \arA23[11] [4], \arA23[11] [3],
       \arA23[11] [2], \arA23[11] [1], 1'b1}), .in_12 ({\arA23[12] [9],
       \arA23[12] [8], \arA23[12] [7], \arA23[12] [6], 1'b0,
       \arA23[12] [4], \arA23[12] [3], \arA23[12] [2], \arA23[12] [1],
       \arA23[12] [0]}), .in_13 ({\arA23[13] [9], \arA23[13] [8], 1'b1,
       \arA23[13] [6], 1'b0, \arA23[13] [4], \arA23[13] [3],
       \arA23[13] [2], \arA23[13] [1], 1'b1}), .in_14 (10'b1111000111),
       .in_15 ({_X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_}), .z
       (plaA2));
  fx68k_mux_1316 \mux_arA1[0]_411_10 (.ctl ({n_23665, n_23666, n_23667,
       n_23668, n_23669, n_23670, n_23671}), .in_0 (5'b00111), .in_1
       (5'b00111), .in_2 (5'b00111), .in_3 (5'b00111), .in_4
       (5'b00111), .in_5 (5'b00111), .in_6 (5'b11000), .z ({n_25163,
       n_25154, n_25145, n_25140, n_25127}));
  fx68k_mux_290 \mux_arA1[0]_339_24 (.ctl ({n_41, n_83, n_125, n_167,
       n_23682}), .in_0 ({n_25164, n_25159, n_25155, n_25150, n_25146,
       n_25141, n_25136, n_25132, n_25128, n_25123}), .in_1 ({n_25165,
       n_25160, n_25156, n_25151, n_25147, n_25142, n_25137, n_25133,
       n_25129, n_25124}), .in_2 ({n_25166, n_25161, n_25157, n_25152,
       n_25148, n_25143, n_25138, n_25134, n_25130, n_25125}), .in_3
       ({n_25167, n_25162, n_25158, n_25153, n_25149, n_25144, n_25139,
       n_25135, n_25131, n_25126}), .in_4 ({1'b1, n_25163, 1'b1,
       n_25154, 1'b1, n_25145, n_25140, 2'b00, n_25127}), .z ({n_25177,
       n_25176, n_25175, n_25174, n_25173, n_25172, n_25171, n_25170,
       n_25169, n_25168}));
  fx68k_mux_290 \mux_arA1[0]_267_24 (.ctl ({n_23697, n_23698, n_23699,
       n_23700, n_23701}), .in_0 (10'b1111100000), .in_1
       (10'b1010111001), .in_2 (10'b1010111001), .in_3
       (10'b1111100000), .in_4 ({n_25177, n_25176, n_25175, n_25174,
       n_25173, n_25172, n_25171, n_25170, n_25169, n_25168}), .z
       ({n_25187, n_25186, n_25185, n_25184, n_25183, n_25182, n_25181,
       n_25180, n_25179, n_25178}));
  fx68k_bmux_299 \mux_arA1[0]_249_32 (.ctl (n_23521), .in_0 ({n_25187,
       n_25186, n_25185, n_25184, n_25183, n_25182, n_25181, n_25180,
       n_25179, n_25178}), .in_1 (10'b1111100000), .z ({n_25197,
       n_25196, n_25195, n_25194, n_25193, n_25192, n_25191, n_25190,
       n_25189, n_25188}));
  fx68k_bmux_299 \mux_arA1[0]_231_32 (.ctl (n_23511), .in_0 ({n_25197,
       n_25196, n_25195, n_25194, n_25193, n_25192, n_25191, n_25190,
       n_25189, n_25188}), .in_1 (10'b1010111001), .z ({n_25207,
       n_25206, n_25205, n_25204, n_25203, n_25202, n_25201, n_25200,
       n_25199, n_25198}));
  fx68k_bmux_299 \mux_arA1[0]_213_32 (.ctl (n_23501), .in_0 ({n_25207,
       n_25206, n_25205, n_25204, n_25203, n_25202, n_25201, n_25200,
       n_25199, n_25198}), .in_1 (10'b1010111001), .z ({n_25217,
       n_25216, n_25215, n_25214, n_25213, n_25212, n_25211, n_25210,
       n_25209, n_25208}));
  fx68k_bmux_299 \mux_arA1[0]_195_32 (.ctl (n_23491), .in_0 ({n_25217,
       n_25216, n_25215, n_25214, n_25213, n_25212, n_25211, n_25210,
       n_25209, n_25208}), .in_1 (10'b1010111001), .z ({n_25227,
       n_25226, n_25225, n_25224, n_25223, n_25222, n_25221, n_25220,
       n_25219, n_25218}));
  fx68k_bmux_299 \mux_arA1[0]_177_27 (.ctl (n_23477), .in_0 ({n_25227,
       n_25226, n_25225, n_25224, n_25223, n_25222, n_25221, n_25220,
       n_25219, n_25218}), .in_1 (10'b1010111001), .z ({\arA1[0] [9],
       \arA1[0] [8], \arA1[0] [7], \arA1[0] [6], \arA1[0] [5],
       \arA1[0] [4], \arA1[0] [3], \arA1[0] [2], \arA1[0] [1],
       \arA1[0] [0]}));
  fx68k_mux_93 \mux_arA1[1]_902_14 (.ctl ({n_24058, n_24059, n_24060,
       n_24061, n_24062, n_24063, n_24064, n_24065}), .in_0
       ({\cmbsop_arA1[1] [19], \cmbsop_arA1[1] [18],
       \cmbsop_arA1[1] [17], \cmbsop_arA1[1] [16], \cmbsop_arA1[1]
       [15], \cmbsop_arA1[1] [14], \cmbsop_arA1[1] [13],
       \cmbsop_arA1[1] [12], \cmbsop_arA1[1] [11], \cmbsop_arA1[1]
       [10]}), .in_1 ({n_25291, n_25284, n_25277, n_25270, n_25263,
       n_25256, n_25249, n_25242, n_25235, n_25228}), .in_2 ({n_25292,
       n_25285, n_25278, n_25271, n_25264, n_25257, n_25250, n_25243,
       n_25236, n_25229}), .in_3 ({n_25293, n_25286, n_25279, n_25272,
       n_25265, n_25258, n_25251, n_25244, n_25237, n_25230}), .in_4
       ({n_25294, n_25287, n_25280, n_25273, n_25266, n_25259, n_25252,
       n_25245, n_25238, n_25231}), .in_5 ({n_25295, n_25288, n_25281,
       n_25274, n_25267, n_25260, n_25253, n_25246, n_25239, n_25232}),
       .in_6 ({n_25296, n_25289, n_25282, n_25275, n_25268, n_25261,
       n_25254, n_25247, n_25240, n_25233}), .in_7 ({n_25297, n_25290,
       n_25283, n_25276, n_25269, n_25262, n_25255, n_25248, n_25241,
       n_25234}), .z ({\arA1[1] [9], \arA1[1] [8], \arA1[1] [7],
       \arA1[1] [6], \arA1[1] [5], \arA1[1] [4], \arA1[1] [3],
       \arA1[1] [2], \arA1[1] [1], \arA1[1] [0]}));
  fx68k_bmux_1352 \mux_arA1[2]_1045_14 (.ctl (movEa), .in_0 ({1'b0,
       \cmbsop_arA1[2] [18], \cmbsop_arA1[2] [17], \cmbsop_arA1[2]
       [16], \cmbsop_arA1[2] [15], \cmbsop_arA1[2] [14],
       \cmbsop_arA1[2] [13], \cmbsop_arA1[2] [12], \cmbsop_arA1[2]
       [11], \cmbsop_arA1[2] [10]}), .in_1 ({1'b0, n_25362, n_25354,
       n_25346, n_25338, n_25330, n_25322, n_25314, n_25306, n_25298}),
       .in_2 ({n_25370, n_25363, n_25355, n_25347, n_25339, n_25331,
       n_25323, n_25315, n_25307, n_25299}), .in_3 ({n_25371, n_25364,
       n_25356, n_25348, n_25340, n_25332, n_25324, n_25316, n_25308,
       n_25300}), .in_4 ({n_25372, n_25365, n_25357, n_25349, n_25341,
       n_25333, n_25325, n_25317, n_25309, n_25301}), .in_5 ({n_25373,
       n_25366, n_25358, n_25350, n_25342, n_25334, n_25326, n_25318,
       n_25310, n_25302}), .in_6 ({1'b0, n_25367, n_25359, n_25351,
       n_25343, n_25335, n_25327, n_25319, n_25311, n_25303}), .in_7
       ({n_25374, n_25368, n_25360, n_25352, n_25344, n_25336, n_25328,
       n_25320, n_25312, n_25304}), .in_8 ({1'b0, n_25369, n_25361,
       n_25353, n_25345, n_25337, n_25329, n_25321, n_25313, n_25305}),
       .z ({\arA1[2] [9], \arA1[2] [8], \arA1[2] [7], \arA1[2] [6],
       \arA1[2] [5], \arA1[2] [4], \arA1[2] [3], \arA1[2] [2],
       \arA1[2] [1], \arA1[2] [0]}));
  fx68k_bmux_1352 \mux_arA1[3]_1205_14 (.ctl (movEa), .in_0
       ({\cmbsop_arA1[3] [19], \cmbsop_arA1[3] [18],
       \cmbsop_arA1[3] [17], \cmbsop_arA1[3] [16], \cmbsop_arA1[3]
       [15], \cmbsop_arA1[3] [14], \cmbsop_arA1[3] [13],
       \cmbsop_arA1[3] [12], \cmbsop_arA1[3] [11], \cmbsop_arA1[3]
       [10]}), .in_1 ({n_25447, n_25439, n_25431, n_25423, n_25415,
       n_25407, n_25399, n_25391, n_25383, n_25375}), .in_2 ({n_25448,
       n_25440, n_25432, n_25424, n_25416, n_25408, n_25400, n_25392,
       n_25384, n_25376}), .in_3 ({n_25449, n_25441, n_25433, n_25425,
       n_25417, n_25409, n_25401, n_25393, n_25385, n_25377}), .in_4
       ({n_25450, n_25442, n_25434, n_25426, n_25418, n_25410, n_25402,
       n_25394, n_25386, n_25378}), .in_5 ({n_25451, n_25443, n_25435,
       n_25427, n_25419, n_25411, n_25403, n_25395, n_25387, n_25379}),
       .in_6 ({n_25452, n_25444, n_25436, n_25428, n_25420, n_25412,
       n_25404, n_25396, n_25388, n_25380}), .in_7 ({n_25453, n_25445,
       n_25437, n_25429, n_25421, n_25413, n_25405, n_25397, n_25389,
       n_25381}), .in_8 ({n_25454, n_25446, n_25438, n_25430, n_25422,
       n_25414, n_25406, n_25398, n_25390, n_25382}), .z ({\arA1[3]
       [9], \arA1[3] [8], \arA1[3] [7], \arA1[3] [6], \arA1[3] [5],
       \arA1[3] [4], \arA1[3] [3], \arA1[3] [2], \arA1[3] [1],
       \arA1[3] [0]}));
  fx68k_case_box_374 ctl_674_19(.in_0 (col), .out_0 ({n_25455,
       UNCONNECTED334, n_25456, UNCONNECTED333, UNCONNECTED332,
       n_25457, n_25458, n_25459, n_25460, n_25461, n_25462,
       UNCONNECTED331, UNCONNECTED330}));
  fx68k_mux_1354 \mux_cmbsop_arA1[4]_674_19 (.ctl ({n_25455, n_25456,
       n_25457, n_25458, n_25459, n_25460, n_25461, n_25462}), .in_0
       (18'b100000010000000000), .in_1 (18'b001111000000000000), .in_2
       (18'b001111010000000000), .in_3 (18'b011111110000000000), .in_4
       (18'b001110000000000000), .in_5 (18'b011110100000000000), .in_6
       (18'b001111010000000000), .in_7 (18'b011111110000000000), .z
       ({n_25698, n_25676, n_25655, n_25643, n_25631, n_25619, n_25607,
       n_25595, UNCONNECTED344, UNCONNECTED343, UNCONNECTED342,
       UNCONNECTED341, UNCONNECTED340, UNCONNECTED339, UNCONNECTED338,
       UNCONNECTED337, UNCONNECTED336, UNCONNECTED335}));
  fx68k_case_box_377 ctl_692_19(.in_0 (col), .out_0 ({n_25463,
       UNCONNECTED350, n_25464, UNCONNECTED349, n_25465, n_25466,
       n_25467, n_25468, n_25469, UNCONNECTED348, UNCONNECTED347,
       UNCONNECTED346, UNCONNECTED345}));
  fx68k_mux_1371 \mux_cmbsop_arA1[4]_692_19 (.ctl ({n_25463, n_25464,
       n_25465, n_25466, n_25467, n_25468, n_25469}), .in_0
       (18'b000100110000000000), .in_1 (18'b110000000000000000), .in_2
       (18'b110001000000000000), .in_3 (18'b011100010000000000), .in_4
       (18'b100001010000000000), .in_5 (18'b011011010000000000), .in_6
       (18'b011001010000000000), .z ({n_25699, n_25677, n_25665,
       n_25644, n_25632, n_25620, n_25608, n_25596, UNCONNECTED360,
       UNCONNECTED359, UNCONNECTED358, UNCONNECTED357, UNCONNECTED356,
       UNCONNECTED355, UNCONNECTED354, UNCONNECTED353, UNCONNECTED352,
       UNCONNECTED351}));
  fx68k_case_box_380 ctl_710_19(.in_0 (col), .out_0 ({n_25470,
       UNCONNECTED366, n_25471, UNCONNECTED365, n_25472, n_25473,
       n_25474, n_25475, n_25476, UNCONNECTED364, UNCONNECTED363,
       UNCONNECTED362, UNCONNECTED361}));
  fx68k_mux_1388 \mux_cmbsop_arA1[4]_710_19 (.ctl ({n_25470, n_25471,
       n_25472, n_25473, n_25474, n_25475, n_25476}), .in_0
       (19'b1000100100000000000), .in_1 (19'b1110000000000000000),
       .in_2 (19'b1110001000000000000), .in_3
       (19'b0111100010000000000), .in_4 (19'b1100001010000000000),
       .in_5 (19'b0111011010000000000), .in_6
       (19'b0111001010000000000), .z ({n_25700, n_25688, n_25678,
       n_25666, n_25645, n_25633, n_25621, n_25609, n_25597,
       UNCONNECTED376, UNCONNECTED375, UNCONNECTED374, UNCONNECTED373,
       UNCONNECTED372, UNCONNECTED371, UNCONNECTED370, UNCONNECTED369,
       UNCONNECTED368, UNCONNECTED367}));
  fx68k_case_box_383 ctl_836_19(.in_0 (col), .out_0 ({UNCONNECTED382,
       UNCONNECTED381, n_25477, UNCONNECTED380, UNCONNECTED379,
       n_25478, n_25479, n_25480, n_25481, n_25482, n_25483,
       UNCONNECTED378, UNCONNECTED377}));
  fx68k_mux_1371 \mux_cmbsop_arA1[4]_836_19 (.ctl ({n_25477, n_25478,
       n_25479, n_25480, n_25481, n_25482, n_25483}), .in_0
       (18'b101100010000000000), .in_1 (18'b101100100000000000), .in_2
       (18'b011110110000000000), .in_3 (18'b100101010000000000), .in_4
       (18'b111001000000000000), .in_5 (18'b101100100000000000), .in_6
       (18'b011110110000000000), .z ({n_25570, n_25567, n_25564,
       n_25557, n_25554, n_25551, n_25548, n_25545, UNCONNECTED392,
       UNCONNECTED391, UNCONNECTED390, UNCONNECTED389, UNCONNECTED388,
       UNCONNECTED387, UNCONNECTED386, UNCONNECTED385, UNCONNECTED384,
       UNCONNECTED383}));
  fx68k_case_box_386 ctl_854_19(.in_0 (col), .out_0 ({UNCONNECTED398,
       UNCONNECTED397, n_25484, UNCONNECTED396, UNCONNECTED395,
       n_25485, n_25486, n_25487, n_25488, n_25489, n_25490,
       UNCONNECTED394, UNCONNECTED393}));
  fx68k_mux_1423 \mux_cmbsop_arA1[4]_854_19 (.ctl ({n_25484, n_25485,
       n_25486, n_25487, n_25488, n_25489, n_25490}), .in_0
       (17'b10011110000000000), .in_1 (17'b10101000000000000), .in_2
       (17'b01111110000000000), .in_3 (17'b10100110000000000), .in_4
       (17'b01111100000000000), .in_5 (17'b10101000000000000), .in_6
       (17'b01111110000000000), .z ({n_25533, n_25531, n_25529,
       n_25527, n_25525, n_25523, n_25521, UNCONNECTED408,
       UNCONNECTED407, UNCONNECTED406, UNCONNECTED405, UNCONNECTED404,
       UNCONNECTED403, UNCONNECTED402, UNCONNECTED401, UNCONNECTED400,
       UNCONNECTED399}));
  fx68k_case_box_389 ctl_872_19(.in_0 (col), .out_0 ({UNCONNECTED414,
       UNCONNECTED413, n_25491, UNCONNECTED412, UNCONNECTED411,
       n_25492, n_25493, n_25494, n_25495, n_25496, n_25497,
       UNCONNECTED410, UNCONNECTED409}));
  fx68k_mux_1423 \mux_cmbsop_arA1[4]_872_19 (.ctl ({n_25491, n_25492,
       n_25493, n_25494, n_25495, n_25496, n_25497}), .in_0
       (17'b10010010000000000), .in_1 (17'b10101000000000000), .in_2
       (17'b01111110000000000), .in_3 (17'b10100110000000000), .in_4
       (17'b01111100000000000), .in_5 (17'b10101000000000000), .in_6
       (17'b01111110000000000), .z ({n_25534, n_25532, n_25530,
       n_25528, n_25526, n_25524, n_25522, UNCONNECTED424,
       UNCONNECTED423, UNCONNECTED422, UNCONNECTED421, UNCONNECTED420,
       UNCONNECTED419, UNCONNECTED418, UNCONNECTED417, UNCONNECTED416,
       UNCONNECTED415}));
  fx68k_case_box_392 ctl_152_16(.in_0 (opcode[2:0]), .out_0 ({n_25501,
       n_25502, n_25503, n_25504, n_25505, n_25506, n_25507, n_25508}));
  fx68k_mux_77 mux_cmbsop_a1Misc_152_16(.ctl ({n_25501, n_25502,
       n_25503, n_25504, n_25505, n_25506, n_25507, n_25508}), .in_0
       (9'b000111010), .in_1 (9'b111001100), .in_2 (9'b110100110),
       .in_3 (9'b111000100), .in_4 (9'b010010100), .in_5
       (9'b010010100), .in_6 (9'b010001100), .in_7 ({_X_, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_, 1'b1}), .z ({cmbsop_a1Misc[10:7],
       cmbsop_a1Misc[4:0]}));
  fx68k_mux_1463 mux_a1Misc_143_13(.ctl ({n_25512, n_25513, n_25514,
       n_25515, n_25516, n_25517}), .in_0 (2'b01), .in_1 (2'b00), .in_2
       (2'b01), .in_3 (2'b11), .in_4 (2'b11), .in_5 (2'b10), .z
       (a1Misc[5:4]));
  fx68k_bmux_1464 mux_a1Misc_143_32(.ctl (opcode[5:3]), .in_0
       (8'b01110000), .in_1 (8'b01110000), .in_2 (8'b11001011), .in_3
       (8'b01001001), .in_4 (8'b10110101), .in_5 (8'b10000000), .in_6
       ({cmbsop_a1Misc[10:7], cmbsop_a1Misc[4:1]}), .z ({a1Misc[9:6],
       a1Misc[3:0]}));
  fx68k_case_box_398 ctl_opcode_853_10(.in_0 (opcode[11:6]), .out_0
       ({n_25518, n_25519, n_25520, n_26717}));
  fx68k_mux_1465 \mux_arA1[4]_853_10 (.ctl ({n_25518, n_25519,
       n_25520}), .in_0 ({n_25533, n_25531, n_25529, n_25527, n_25525,
       3'b100, n_25523, n_25521}), .in_1 ({n_25534, n_25532, n_25530,
       n_25528, n_25526, 3'b101, n_25524, n_25522}), .in_2 (a1Misc), .z
       ({n_25571, n_25568, n_25565, n_25562, n_25560, n_25558, n_25555,
       n_25552, n_25549, n_25546}));
  fx68k_mux_1465 \mux_arA1[4]_817_24 (.ctl ({n_167, n_125, n_25543}),
       .in_0 ({n_25569, n_25566, n_25563, n_25561, n_25559, n_25556,
       n_25553, n_25550, n_25547, n_25544}), .in_1 ({n_25570, n_25567,
       n_25564, 2'b11, n_25557, n_25554, n_25551, n_25548, n_25545}),
       .in_2 ({n_25571, n_25568, n_25565, n_25562, n_25560, n_25558,
       n_25555, n_25552, n_25549, n_25546}), .z ({n_25587, n_25586,
       n_25585, n_25583, n_25581, n_25580, n_25578, n_25576, n_25574,
       n_25572}));
  fx68k_bmux_299 \mux_arA1[4]_799_32 (.ctl (n_24491), .in_0 ({n_25587,
       n_25586, n_25585, n_25583, n_25581, n_25580, n_25578, n_25576,
       n_25574, n_25572}), .in_1 ({2'b01, n_25584, n_25582, 1'b1,
       n_25579, n_25577, n_25575, n_25573, 1'b1}), .z ({n_25704,
       n_25693, n_25683, n_25671, n_25660, n_25650, n_25638, n_25626,
       n_25614, n_25602}));
  fx68k_mux_119 \mux_arA1[4]_601_10 (.ctl ({n_24511, n_24512, n_24513,
       n_24514, n_25588, n_25589, n_25590, n_24515, n_24516, n_24517,
       n_24518, n_24519}), .in_0 ({n_25694, n_25684, n_25672, n_25661,
       n_25651, n_25639, n_25627, n_25615, n_25603, n_25591}), .in_1
       ({n_25695, n_25685, n_25673, n_25662, n_25652, n_25640, n_25628,
       n_25616, n_25604, n_25592}), .in_2 ({n_25696, n_25686, n_25674,
       n_25663, n_25653, n_25641, n_25629, n_25617, n_25605, n_25593}),
       .in_3 ({n_25697, n_25687, n_25675, n_25664, n_25654, n_25642,
       n_25630, n_25618, n_25606, n_25594}), .in_4 ({n_25698, 1'b1,
       n_25676, 1'b1, n_25655, n_25643, n_25631, n_25619, n_25607,
       n_25595}), .in_5 ({n_25699, 1'b1, n_25677, n_25665, 1'b1,
       n_25644, n_25632, n_25620, n_25608, n_25596}), .in_6 ({n_25700,
       n_25688, n_25678, n_25666, 1'b1, n_25645, n_25633, n_25621,
       n_25609, n_25597}), .in_7 ({n_25701, n_25689, n_25679, n_25667,
       n_25656, n_25646, n_25634, n_25622, n_25610, n_25598}), .in_8
       ({n_25702, n_25690, n_25680, n_25668, n_25657, n_25647, n_25635,
       n_25623, n_25611, n_25599}), .in_9 ({1'b0, n_25691, n_25681,
       n_25669, n_25658, n_25648, n_25636, n_25624, n_25612, n_25600}),
       .in_10 ({n_25703, n_25692, n_25682, n_25670, n_25659, n_25649,
       n_25637, n_25625, n_25613, n_25601}), .in_11 ({n_25704, n_25693,
       n_25683, n_25671, n_25660, n_25650, n_25638, n_25626, n_25614,
       n_25602}), .z ({n_25733, n_25731, n_25728, n_25725, n_25722,
       n_25719, n_25716, n_25713, n_25710, n_25707}));
  fx68k_mux_812 \mux_arA1[4]_547_19 (.ctl ({n_24536, n_24537, n_24538,
       n_24539}), .in_0 ({\cmbsop_arA1[4] [19], \cmbsop_arA1[4] [18],
       \cmbsop_arA1[4] [17], \cmbsop_arA1[4] [16], \cmbsop_arA1[4]
       [15], \cmbsop_arA1[4] [14], \cmbsop_arA1[4] [13],
       \cmbsop_arA1[4] [12], \cmbsop_arA1[4] [11], \cmbsop_arA1[4]
       [10]}), .in_1 ({n_25732, n_25729, n_25726, n_25723, n_25720,
       n_25717, n_25714, n_25711, n_25708, n_25705}), .in_2 ({1'b0,
       n_25730, n_25727, n_25724, n_25721, n_25718, n_25715, n_25712,
       n_25709, n_25706}), .in_3 ({n_25733, n_25731, n_25728, n_25725,
       n_25722, n_25719, n_25716, n_25713, n_25710, n_25707}), .z
       ({\arA1[4] [9], \arA1[4] [8], \arA1[4] [7], \arA1[4] [6],
       \arA1[4] [5], \arA1[4] [4], \arA1[4] [3], \arA1[4] [2],
       \arA1[4] [1], \arA1[4] [0]}));
  fx68k_bmux_1502 \mux_arA1[5]_1365_14 (.ctl (opcode[8:6]), .in_0
       ({\cmbsop_arA1[5] [19], \cmbsop_arA1[5] [18],
       \cmbsop_arA1[5] [17], \cmbsop_arA1[5] [16], \cmbsop_arA1[5]
       [15], \cmbsop_arA1[5] [14], \cmbsop_arA1[5] [13],
       \cmbsop_arA1[5] [12], \cmbsop_arA1[5] [11], \cmbsop_arA1[5]
       [10]}), .in_1 ({n_25797, n_25790, n_25783, n_25776, n_25769,
       n_25762, n_25755, n_25748, n_25741, n_25734}), .in_2 ({n_25798,
       n_25791, n_25784, n_25777, n_25770, n_25763, n_25756, n_25749,
       n_25742, n_25735}), .in_3 ({n_25799, n_25792, n_25785, n_25778,
       n_25771, n_25764, n_25757, n_25750, n_25743, n_25736}), .in_4
       ({n_25800, n_25793, n_25786, n_25779, n_25772, n_25765, n_25758,
       n_25751, n_25744, n_25737}), .in_5 ({n_25801, n_25794, n_25787,
       n_25780, n_25773, n_25766, n_25759, n_25752, n_25745, n_25738}),
       .in_6 ({n_25802, n_25795, n_25788, n_25781, n_25774, n_25767,
       n_25760, n_25753, n_25746, n_25739}), .in_7 ({n_25803, n_25796,
       n_25789, n_25782, n_25775, n_25768, n_25761, n_25754, n_25747,
       n_25740}), .z ({\arA1[5] [9], \arA1[5] [8], \arA1[5] [7],
       \arA1[5] [6], \arA1[5] [5], \arA1[5] [4], \arA1[5] [3],
       \arA1[5] [2], \arA1[5] [1], \arA1[5] [0]}));
  fx68k_bmux_1503 mux_88_24(.ctl (n_25805), .in_0 (1'b1), .in_1 (1'b0),
       .z (n_25807));
  fx68k_bmux_1504 mux_90_24(.ctl (n_25806), .in_0 (4'b0011), .in_1
       (4'b1100), .z ({n_25811, n_25810, n_25809, n_25808}));
  fx68k_bmux_1505 \mux_arA1[6]_87_25 (.ctl (n_25804), .in_0 ({n_25811,
       n_25810, 1'b0, n_25809, n_25808, 1'b0}), .in_1 ({4'b0010,
       n_25807, 1'b1}), .z ({\arA1[6] [9], \arA1[6] [8], \arA1[6] [7],
       \arA1[6] [6], \arA1[6] [5], \arA1[6] [0]}));
  fx68k_bmux_1502 \mux_arA1[8]_1483_14 (.ctl (opcode[8:6]), .in_0
       ({\cmbsop_arA1[8] [19], \cmbsop_arA1[8] [18],
       \cmbsop_arA1[8] [17], \cmbsop_arA1[8] [16], \cmbsop_arA1[8]
       [15], \cmbsop_arA1[8] [14], \cmbsop_arA1[8] [13],
       \cmbsop_arA1[8] [12], \cmbsop_arA1[8] [11], \cmbsop_arA1[8]
       [10]}), .in_1 ({n_25875, n_25868, n_25861, n_25854, n_25847,
       n_25840, n_25833, n_25826, n_25819, n_25812}), .in_2 ({1'b0,
       n_25869, n_25862, n_25855, n_25848, n_25841, n_25834, n_25827,
       n_25820, n_25813}), .in_3 ({n_25876, n_25870, n_25863, n_25856,
       n_25849, n_25842, n_25835, n_25828, n_25821, n_25814}), .in_4
       ({n_25877, n_25871, n_25864, n_25857, n_25850, n_25843, n_25836,
       n_25829, n_25822, n_25815}), .in_5 ({n_25878, n_25872, n_25865,
       n_25858, n_25851, n_25844, n_25837, n_25830, n_25823, n_25816}),
       .in_6 ({1'b0, n_25873, n_25866, n_25859, n_25852, n_25845,
       n_25838, n_25831, n_25824, n_25817}), .in_7 ({n_25879, n_25874,
       n_25867, n_25860, n_25853, n_25846, n_25839, n_25832, n_25825,
       n_25818}), .z ({\arA1[8] [9], \arA1[8] [8], \arA1[8] [7],
       \arA1[8] [6], \arA1[8] [5], \arA1[8] [4], \arA1[8] [3],
       \arA1[8] [2], \arA1[8] [1], \arA1[8] [0]}));
  fx68k_bmux_1502 \mux_arA1[9]_1625_14 (.ctl (opcode[8:6]), .in_0
       ({\cmbsop_arA1[9] [19], \cmbsop_arA1[9] [18],
       \cmbsop_arA1[9] [17], \cmbsop_arA1[9] [16], \cmbsop_arA1[9]
       [15], \cmbsop_arA1[9] [14], \cmbsop_arA1[9] [13],
       \cmbsop_arA1[9] [12], \cmbsop_arA1[9] [11], \cmbsop_arA1[9]
       [10]}), .in_1 ({n_25943, n_25936, n_25929, n_25922, n_25915,
       n_25908, n_25901, n_25894, n_25887, n_25880}), .in_2 ({1'b0,
       n_25937, n_25930, n_25923, n_25916, n_25909, n_25902, n_25895,
       n_25888, n_25881}), .in_3 ({n_25944, n_25938, n_25931, n_25924,
       n_25917, n_25910, n_25903, n_25896, n_25889, n_25882}), .in_4
       ({n_25945, n_25939, n_25932, n_25925, n_25918, n_25911, n_25904,
       n_25897, n_25890, n_25883}), .in_5 ({n_25946, n_25940, n_25933,
       n_25926, n_25919, n_25912, n_25905, n_25898, n_25891, n_25884}),
       .in_6 ({1'b0, n_25941, n_25934, n_25927, n_25920, n_25913,
       n_25906, n_25899, n_25892, n_25885}), .in_7 ({1'b0, n_25942,
       n_25935, n_25928, n_25921, n_25914, n_25907, n_25900, n_25893,
       n_25886}), .z ({\arA1[9] [9], \arA1[9] [8], \arA1[9] [7],
       \arA1[9] [6], \arA1[9] [5], \arA1[9] [4], \arA1[9] [3],
       \arA1[9] [2], \arA1[9] [1], \arA1[9] [0]}));
  fx68k_bmux_1502 \mux_arA1[11]_1767_14 (.ctl (opcode[8:6]), .in_0
       ({\cmbsop_arA1[11] [19], \cmbsop_arA1[11] [18],
       \cmbsop_arA1[11] [17], \cmbsop_arA1[11] [16],
       \cmbsop_arA1[11] [15], \cmbsop_arA1[11] [14],
       \cmbsop_arA1[11] [13], \cmbsop_arA1[11] [12],
       \cmbsop_arA1[11] [11], \cmbsop_arA1[11] [10]}), .in_1 ({n_26010,
       n_26003, n_25996, n_25989, n_25982, n_25975, n_25968, n_25961,
       n_25954, n_25947}), .in_2 ({1'b0, n_26004, n_25997, n_25990,
       n_25983, n_25976, n_25969, n_25962, n_25955, n_25948}), .in_3
       ({n_26011, n_26005, n_25998, n_25991, n_25984, n_25977, n_25970,
       n_25963, n_25956, n_25949}), .in_4 ({n_26012, n_26006, n_25999,
       n_25992, n_25985, n_25978, n_25971, n_25964, n_25957, n_25950}),
       .in_5 ({n_26013, n_26007, n_26000, n_25993, n_25986, n_25979,
       n_25972, n_25965, n_25958, n_25951}), .in_6 ({1'b0, n_26008,
       n_26001, n_25994, n_25987, n_25980, n_25973, n_25966, n_25959,
       n_25952}), .in_7 ({1'b0, n_26009, n_26002, n_25995, n_25988,
       n_25981, n_25974, n_25967, n_25960, n_25953}), .z ({\arA1[11]
       [9], \arA1[11] [8], \arA1[11] [7], \arA1[11] [6], \arA1[11] [5],
       \arA1[11] [4], \arA1[11] [3], \arA1[11] [2], \arA1[11] [1],
       \arA1[11] [0]}));
  fx68k_bmux_1502 \mux_arA1[12]_1909_14 (.ctl (opcode[8:6]), .in_0
       ({\cmbsop_arA1[12] [19], \cmbsop_arA1[12] [18],
       \cmbsop_arA1[12] [17], \cmbsop_arA1[12] [16],
       \cmbsop_arA1[12] [15], \cmbsop_arA1[12] [14],
       \cmbsop_arA1[12] [13], \cmbsop_arA1[12] [12],
       \cmbsop_arA1[12] [11], \cmbsop_arA1[12] [10]}), .in_1 ({n_26077,
       n_26070, n_26063, n_26056, n_26049, n_26042, n_26035, n_26028,
       n_26021, n_26014}), .in_2 ({1'b0, n_26071, n_26064, n_26057,
       n_26050, n_26043, n_26036, n_26029, n_26022, n_26015}), .in_3
       ({n_26078, n_26072, n_26065, n_26058, n_26051, n_26044, n_26037,
       n_26030, n_26023, n_26016}), .in_4 ({n_26079, n_26073, n_26066,
       n_26059, n_26052, n_26045, n_26038, n_26031, n_26024, n_26017}),
       .in_5 ({n_26080, n_26074, n_26067, n_26060, n_26053, n_26046,
       n_26039, n_26032, n_26025, n_26018}), .in_6 ({n_26081, n_26075,
       n_26068, n_26061, n_26054, n_26047, n_26040, n_26033, n_26026,
       n_26019}), .in_7 ({n_26082, n_26076, n_26069, n_26062, n_26055,
       n_26048, n_26041, n_26034, n_26027, n_26020}), .z ({\arA1[12]
       [9], \arA1[12] [8], \arA1[12] [7], \arA1[12] [6], \arA1[12] [5],
       \arA1[12] [4], \arA1[12] [3], \arA1[12] [2], \arA1[12] [1],
       \arA1[12] [0]}));
  fx68k_bmux_1502 \mux_arA1[13]_2051_14 (.ctl (opcode[8:6]), .in_0
       ({\cmbsop_arA1[13] [19], \cmbsop_arA1[13] [18],
       \cmbsop_arA1[13] [17], \cmbsop_arA1[13] [16],
       \cmbsop_arA1[13] [15], \cmbsop_arA1[13] [14],
       \cmbsop_arA1[13] [13], \cmbsop_arA1[13] [12],
       \cmbsop_arA1[13] [11], \cmbsop_arA1[13] [10]}), .in_1 ({n_26146,
       n_26139, n_26132, n_26125, n_26118, n_26111, n_26104, n_26097,
       n_26090, n_26083}), .in_2 ({1'b0, n_26140, n_26133, n_26126,
       n_26119, n_26112, n_26105, n_26098, n_26091, n_26084}), .in_3
       ({n_26147, n_26141, n_26134, n_26127, n_26120, n_26113, n_26106,
       n_26099, n_26092, n_26085}), .in_4 ({n_26148, n_26142, n_26135,
       n_26128, n_26121, n_26114, n_26107, n_26100, n_26093, n_26086}),
       .in_5 ({n_26149, n_26143, n_26136, n_26129, n_26122, n_26115,
       n_26108, n_26101, n_26094, n_26087}), .in_6 ({1'b0, n_26144,
       n_26137, n_26130, n_26123, n_26116, n_26109, n_26102, n_26095,
       n_26088}), .in_7 ({1'b0, n_26145, n_26138, n_26131, n_26124,
       n_26117, n_26110, n_26103, n_26096, n_26089}), .z ({\arA1[13]
       [9], \arA1[13] [8], \arA1[13] [7], \arA1[13] [6], \arA1[13] [5],
       \arA1[13] [4], \arA1[13] [3], \arA1[13] [2], \arA1[13] [1],
       \arA1[13] [0]}));
  fx68k_case_box_404 ctl_col_111_23(.in_0 (col), .out_0 ({n_26150,
       n_26151, n_26152, n_26153, n_26154, n_26155, n_26156, n_26176}));
  fx68k_mux_272 \mux_arA1[14]_111_23 (.ctl ({n_26150, n_26151, n_26152,
       n_26153, n_26154, n_26155, n_26156}), .in_0 (10'b0000000110),
       .in_1 (10'b1000011100), .in_2 (10'b0100000011), .in_3
       (10'b0111000010), .in_4 (10'b0111100011), .in_5
       (10'b0000001010), .in_6 (10'b0111100010), .z ({n_26175, n_26174,
       n_26173, n_26172, n_26171, n_26170, n_26169, n_26167, n_26165,
       n_26163}));
  fx68k_bmux_1520 mux_129_33(.ctl (opcode[5]), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_26161, n_26159}));
  fx68k_bmux_1520 mux_133_33(.ctl (opcode[5]), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_26162, n_26160}));
  fx68k_mux_1522 \mux_arA1[14]_125_23 (.ctl ({n_73, n_26158}), .in_0
       ({1'b0, n_26161, n_26159}), .in_1 ({1'b1, n_26162, n_26160}), .z
       ({n_26168, n_26166, n_26164}));
  fx68k_bmux_299 \mux_arA1[14]_108_35 (.ctl (n_25122), .in_0
       ({7'b1110000, n_26168, n_26166, n_26164}), .in_1 ({n_26175,
       n_26174, n_26173, n_26172, n_26171, n_26170, n_26169, n_26167,
       n_26165, n_26163}), .z ({\arA1[14] [9], \arA1[14] [8],
       \arA1[14] [7], \arA1[14] [6], \arA1[14] [5], \arA1[14] [4],
       \arA1[14] [3], \arA1[14] [2], \arA1[14] [1], \arA1[14] [0]}));
  fx68k_bmux_1313 \mux_arA1[line]_77_19 (.ctl (opcode[15:12]), .in_0
       ({\arA1[0] [9], \arA1[0] [8], \arA1[0] [7], \arA1[0] [6],
       \arA1[0] [5], \arA1[0] [4], \arA1[0] [3], \arA1[0] [2],
       \arA1[0] [1], \arA1[0] [0]}), .in_1 ({\arA1[1] [9], \arA1[1]
       [8], \arA1[1] [7], \arA1[1] [6], \arA1[1] [5], \arA1[1] [4],
       \arA1[1] [3], \arA1[1] [2], \arA1[1] [1], \arA1[1] [0]}), .in_2
       ({\arA1[2] [9], \arA1[2] [8], \arA1[2] [7], \arA1[2] [6],
       \arA1[2] [5], \arA1[2] [4], \arA1[2] [3], \arA1[2] [2],
       \arA1[2] [1], \arA1[2] [0]}), .in_3 ({\arA1[3] [9], \arA1[3]
       [8], \arA1[3] [7], \arA1[3] [6], \arA1[3] [5], \arA1[3] [4],
       \arA1[3] [3], \arA1[3] [2], \arA1[3] [1], \arA1[3] [0]}), .in_4
       ({\arA1[4] [9], \arA1[4] [8], \arA1[4] [7], \arA1[4] [6],
       \arA1[4] [5], \arA1[4] [4], \arA1[4] [3], \arA1[4] [2],
       \arA1[4] [1], \arA1[4] [0]}), .in_5 ({\arA1[5] [9], \arA1[5]
       [8], \arA1[5] [7], \arA1[5] [6], \arA1[5] [5], \arA1[5] [4],
       \arA1[5] [3], \arA1[5] [2], \arA1[5] [1], \arA1[5] [0]}), .in_6
       ({\arA1[6] [9], \arA1[6] [8], \arA1[6] [7], \arA1[6] [6],
       \arA1[6] [5], 4'b0100, \arA1[6] [0]}), .in_7 (10'b1000111011),
       .in_8 ({\arA1[8] [9], \arA1[8] [8], \arA1[8] [7], \arA1[8] [6],
       \arA1[8] [5], \arA1[8] [4], \arA1[8] [3], \arA1[8] [2],
       \arA1[8] [1], \arA1[8] [0]}), .in_9 ({\arA1[9] [9], \arA1[9]
       [8], \arA1[9] [7], \arA1[9] [6], \arA1[9] [5], \arA1[9] [4],
       \arA1[9] [3], \arA1[9] [2], \arA1[9] [1], \arA1[9] [0]}), .in_10
       ({_X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_}), .in_11
       ({\arA1[11] [9], \arA1[11] [8], \arA1[11] [7], \arA1[11] [6],
       \arA1[11] [5], \arA1[11] [4], \arA1[11] [3], \arA1[11] [2],
       \arA1[11] [1], \arA1[11] [0]}), .in_12 ({\arA1[12] [9],
       \arA1[12] [8], \arA1[12] [7], \arA1[12] [6], \arA1[12] [5],
       \arA1[12] [4], \arA1[12] [3], \arA1[12] [2], \arA1[12] [1],
       \arA1[12] [0]}), .in_13 ({\arA1[13] [9], \arA1[13] [8],
       \arA1[13] [7], \arA1[13] [6], \arA1[13] [5], \arA1[13] [4],
       \arA1[13] [3], \arA1[13] [2], \arA1[13] [1], \arA1[13] [0]}),
       .in_14 ({\arA1[14] [9], \arA1[14] [8], \arA1[14] [7],
       \arA1[14] [6], \arA1[14] [5], \arA1[14] [4], \arA1[14] [3],
       \arA1[14] [2], \arA1[14] [1], \arA1[14] [0]}), .in_15 ({_X_,
       _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_}), .z (plaA1));
  fx68k_mux_1526 mux_arIll_111_23(.ctl ({n_26150, n_26151, n_26152,
       n_26153, n_26154, n_26155, n_26156, n_26176}), .in_0 (1'b0),
       .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5
       (1'b0), .in_6 (1'b0), .in_7 (1'b1), .z (n_26178));
  fx68k_mux_1527 mux_arIll_125_23(.ctl ({n_73, n_26158, n_26177}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b1), .z (n_26179));
  fx68k_bmux_1503 mux_arIll_108_35(.ctl (n_25122), .in_0 (n_26179),
       .in_1 (n_26178), .z (arIll[14]));
  fx68k_mux_1529 mux_arIll_178_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26466));
  fx68k_mux_1529 mux_arIll_196_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26464));
  fx68k_mux_1529 mux_arIll_214_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26462));
  fx68k_mux_1529 mux_arIll_232_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26460));
  fx68k_mux_1529 mux_arIll_250_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26458));
  fx68k_mux_1529 mux_arIll_268_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26453));
  fx68k_mux_1529 mux_arIll_286_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26454));
  fx68k_mux_1529 mux_arIll_304_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26455));
  fx68k_mux_1529 mux_arIll_322_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26456));
  fx68k_mux_1529 mux_arIll_340_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26448));
  fx68k_mux_1529 mux_arIll_358_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26449));
  fx68k_mux_1529 mux_arIll_376_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26450));
  fx68k_mux_1529 mux_arIll_394_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26451));
  fx68k_mux_1529 mux_arIll_412_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26441));
  fx68k_mux_1529 mux_arIll_430_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26442));
  fx68k_mux_1529 mux_arIll_448_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26443));
  fx68k_mux_1529 mux_arIll_466_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26444));
  fx68k_mux_1529 mux_arIll_484_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26445));
  fx68k_mux_1529 mux_arIll_502_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26446));
  fx68k_mux_1529 mux_arIll_520_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26447));
  fx68k_mux_1526 mux_arIll_411_10(.ctl ({n_23665, n_23666, n_23667,
       n_23668, n_23669, n_23670, n_23671, n_26440}), .in_0 (n_26441),
       .in_1 (n_26442), .in_2 (n_26443), .in_3 (n_26444), .in_4
       (n_26445), .in_5 (n_26446), .in_6 (n_26447), .in_7 (1'b1), .z
       (n_26452));
  fx68k_mux_1550 mux_arIll_339_24(.ctl ({n_41, n_83, n_125, n_167,
       n_23682}), .in_0 (n_26448), .in_1 (n_26449), .in_2 (n_26450),
       .in_3 (n_26451), .in_4 (n_26452), .z (n_26457));
  fx68k_mux_1550 mux_arIll_267_24(.ctl ({n_23697, n_23698, n_23699,
       n_23700, n_23701}), .in_0 (n_26453), .in_1 (n_26454), .in_2
       (n_26455), .in_3 (n_26456), .in_4 (n_26457), .z (n_26459));
  fx68k_bmux_1503 mux_arIll_249_32(.ctl (n_23521), .in_0 (n_26459),
       .in_1 (n_26458), .z (n_26461));
  fx68k_bmux_1503 mux_arIll_231_32(.ctl (n_23511), .in_0 (n_26461),
       .in_1 (n_26460), .z (n_26463));
  fx68k_bmux_1503 mux_arIll_213_32(.ctl (n_23501), .in_0 (n_26463),
       .in_1 (n_26462), .z (n_26465));
  fx68k_bmux_1503 mux_arIll_195_32(.ctl (n_23491), .in_0 (n_26465),
       .in_1 (n_26464), .z (n_26467));
  fx68k_bmux_1503 mux_arIll_177_27(.ctl (n_23477), .in_0 (n_26467),
       .in_1 (n_26466), .z (arIll[0]));
  fx68k_mux_1529 mux_arIll_548_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26737));
  fx68k_mux_1529 mux_arIll_566_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26738));
  fx68k_mux_1529 mux_arIll_584_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26739));
  fx68k_mux_1529 mux_arIll_602_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26725));
  fx68k_mux_1529 mux_arIll_620_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26726));
  fx68k_mux_1529 mux_arIll_638_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26727));
  fx68k_mux_1529 mux_arIll_656_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26728));
  fx68k_mux_1529 mux_arIll_674_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b1), .in_4 (1'b1), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26729));
  fx68k_mux_1529 mux_arIll_692_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b1), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26730));
  fx68k_mux_1529 mux_arIll_710_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b1), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26731));
  fx68k_mux_1529 mux_arIll_728_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26732));
  fx68k_mux_1529 mux_arIll_746_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26733));
  fx68k_mux_1529 mux_arIll_764_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26734));
  fx68k_mux_1529 mux_arIll_782_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26735));
  fx68k_mux_1529 mux_arIll_800_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b1), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b1), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26723));
  fx68k_mux_1529 mux_arIll_818_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26720));
  fx68k_mux_1529 mux_arIll_836_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b1), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b1), .in_4 (1'b1), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26721));
  fx68k_mux_1529 mux_arIll_854_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b1), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b1), .in_4 (1'b1), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26718));
  fx68k_mux_1529 mux_arIll_872_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b1), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b1), .in_4 (1'b1), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b1), .in_12 (1'b1), .z (n_26719));
  fx68k_mux_1527 mux_illMisc_143_13(.ctl ({n_26715, n_25517, n_26716}),
       .in_0 (1'b0), .in_1 (cmbsop_a1Misc[0]), .in_2 (1'b1), .z
       (illMisc));
  fx68k_mux_1577 mux_arIll_853_10(.ctl ({n_25518, n_25519, n_25520,
       n_26717}), .in_0 (n_26718), .in_1 (n_26719), .in_2 (illMisc),
       .in_3 (1'b1), .z (n_26722));
  fx68k_mux_1527 mux_arIll_817_24(.ctl ({n_167, n_125, n_25543}), .in_0
       (n_26720), .in_1 (n_26721), .in_2 (n_26722), .z (n_26724));
  fx68k_bmux_1503 mux_arIll_799_32(.ctl (n_24491), .in_0 (n_26724),
       .in_1 (n_26723), .z (n_26736));
  fx68k_mux_1580 mux_arIll_601_10(.ctl ({n_24511, n_24512, n_24513,
       n_24514, n_25588, n_25589, n_25590, n_24515, n_24516, n_24517,
       n_24518, n_24519}), .in_0 (n_26725), .in_1 (n_26726), .in_2
       (n_26727), .in_3 (n_26728), .in_4 (n_26729), .in_5 (n_26730),
       .in_6 (n_26731), .in_7 (n_26732), .in_8 (n_26733), .in_9
       (n_26734), .in_10 (n_26735), .in_11 (n_26736), .z (n_26740));
  fx68k_mux_1577 mux_arIll_547_19(.ctl ({n_24536, n_24537, n_24538,
       n_24539}), .in_0 (n_26737), .in_1 (n_26738), .in_2 (n_26739),
       .in_3 (n_26740), .z (arIll[4]));
  fx68k_mux_1529 mux_arIll_905_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26845));
  fx68k_mux_1529 mux_arIll_922_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26846));
  fx68k_mux_1529 mux_arIll_939_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26847));
  fx68k_mux_1529 mux_arIll_956_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26848));
  fx68k_mux_1529 mux_arIll_973_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26849));
  fx68k_mux_1529 mux_arIll_990_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26850));
  fx68k_mux_1529 mux_arIll_1007_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26851));
  fx68k_mux_1529 mux_arIll_1024_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26852));
  fx68k_bmux_1590 mux_arIll_902_14(.ctl (movEa), .in_0 (n_26845), .in_1
       (1'b1), .in_2 (n_26846), .in_3 (n_26847), .in_4 (n_26848), .in_5
       (n_26849), .in_6 (n_26850), .in_7 (n_26851), .in_8 (n_26852),
       .in_9 (1'b1), .in_10 (1'b1), .in_11 (1'b1), .in_12 (1'b1),
       .in_13 (1'b1), .in_14 (1'b1), .in_15 (1'b1), .z (arIll[1]));
  fx68k_mux_1529 mux_arIll_1048_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26970));
  fx68k_mux_1529 mux_arIll_1065_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26971));
  fx68k_mux_1529 mux_arIll_1082_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26972));
  fx68k_mux_1529 mux_arIll_1099_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26973));
  fx68k_mux_1529 mux_arIll_1116_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26974));
  fx68k_mux_1529 mux_arIll_1133_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26975));
  fx68k_mux_1529 mux_arIll_1150_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26976));
  fx68k_mux_1529 mux_arIll_1167_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26977));
  fx68k_mux_1529 mux_arIll_1184_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_26978));
  fx68k_bmux_1590 mux_arIll_1045_14(.ctl (movEa), .in_0 (n_26970),
       .in_1 (n_26971), .in_2 (n_26972), .in_3 (n_26973), .in_4
       (n_26974), .in_5 (n_26975), .in_6 (n_26976), .in_7 (n_26977),
       .in_8 (n_26978), .in_9 (1'b1), .in_10 (1'b1), .in_11 (1'b1),
       .in_12 (1'b1), .in_13 (1'b1), .in_14 (1'b1), .in_15 (1'b1), .z
       (arIll[2]));
  fx68k_mux_1529 mux_arIll_1208_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27096));
  fx68k_mux_1529 mux_arIll_1225_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27097));
  fx68k_mux_1529 mux_arIll_1242_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27098));
  fx68k_mux_1529 mux_arIll_1259_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27099));
  fx68k_mux_1529 mux_arIll_1276_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27100));
  fx68k_mux_1529 mux_arIll_1293_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27101));
  fx68k_mux_1529 mux_arIll_1310_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27102));
  fx68k_mux_1529 mux_arIll_1327_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27103));
  fx68k_mux_1529 mux_arIll_1344_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27104));
  fx68k_bmux_1590 mux_arIll_1205_14(.ctl (movEa), .in_0 (n_27096),
       .in_1 (n_27097), .in_2 (n_27098), .in_3 (n_27099), .in_4
       (n_27100), .in_5 (n_27101), .in_6 (n_27102), .in_7 (n_27103),
       .in_8 (n_27104), .in_9 (1'b1), .in_10 (1'b1), .in_11 (1'b1),
       .in_12 (1'b1), .in_13 (1'b1), .in_14 (1'b1), .in_15 (1'b1), .z
       (arIll[3]));
  fx68k_mux_1611 mux_arIll_1368_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b1), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27185));
  fx68k_mux_1611 mux_arIll_1382_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27186));
  fx68k_mux_1611 mux_arIll_1396_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27187));
  fx68k_mux_1611 mux_arIll_1410_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27188));
  fx68k_mux_1611 mux_arIll_1424_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b1), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27189));
  fx68k_mux_1611 mux_arIll_1438_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27190));
  fx68k_mux_1611 mux_arIll_1452_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27191));
  fx68k_mux_1611 mux_arIll_1466_19(.ctl ({n_27105, n_27106, n_27107,
       n_27108, n_27109, n_27110, n_27111, n_27112, n_27113, n_27114}),
       .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4
       (1'b0), .in_5 (1'b0), .in_6 (1'b0), .in_7 (1'b0), .in_8 (1'b0),
       .in_9 (1'b1), .z (n_27192));
  fx68k_bmux_1619 mux_arIll_1365_14(.ctl (opcode[8:6]), .in_0
       (n_27185), .in_1 (n_27186), .in_2 (n_27187), .in_3 (n_27188),
       .in_4 (n_27189), .in_5 (n_27190), .in_6 (n_27191), .in_7
       (n_27192), .z (arIll[5]));
  fx68k_mux_1529 mux_arIll_1486_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27297));
  fx68k_mux_1529 mux_arIll_1503_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27298));
  fx68k_mux_1529 mux_arIll_1520_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27299));
  fx68k_mux_1529 mux_arIll_1537_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27300));
  fx68k_mux_1529 mux_arIll_1554_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27301));
  fx68k_mux_1529 mux_arIll_1571_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b1), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27302));
  fx68k_mux_1529 mux_arIll_1588_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b1), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27303));
  fx68k_mux_1529 mux_arIll_1605_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27304));
  fx68k_bmux_1619 mux_arIll_1483_14(.ctl (opcode[8:6]), .in_0
       (n_27297), .in_1 (n_27298), .in_2 (n_27299), .in_3 (n_27300),
       .in_4 (n_27301), .in_5 (n_27302), .in_6 (n_27303), .in_7
       (n_27304), .z (arIll[8]));
  fx68k_mux_1529 mux_arIll_1628_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27409));
  fx68k_mux_1529 mux_arIll_1645_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27410));
  fx68k_mux_1529 mux_arIll_1662_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27411));
  fx68k_mux_1529 mux_arIll_1679_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27412));
  fx68k_mux_1529 mux_arIll_1696_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27413));
  fx68k_mux_1529 mux_arIll_1713_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27414));
  fx68k_mux_1529 mux_arIll_1730_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27415));
  fx68k_mux_1529 mux_arIll_1747_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27416));
  fx68k_bmux_1619 mux_arIll_1625_14(.ctl (opcode[8:6]), .in_0
       (n_27409), .in_1 (n_27410), .in_2 (n_27411), .in_3 (n_27412),
       .in_4 (n_27413), .in_5 (n_27414), .in_6 (n_27415), .in_7
       (n_27416), .z (arIll[9]));
  fx68k_mux_1529 mux_arIll_1770_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27521));
  fx68k_mux_1529 mux_arIll_1787_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27522));
  fx68k_mux_1529 mux_arIll_1804_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27523));
  fx68k_mux_1529 mux_arIll_1821_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27524));
  fx68k_mux_1529 mux_arIll_1838_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27525));
  fx68k_mux_1529 mux_arIll_1855_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27526));
  fx68k_mux_1529 mux_arIll_1872_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27527));
  fx68k_mux_1529 mux_arIll_1889_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27528));
  fx68k_bmux_1619 mux_arIll_1767_14(.ctl (opcode[8:6]), .in_0
       (n_27521), .in_1 (n_27522), .in_2 (n_27523), .in_3 (n_27524),
       .in_4 (n_27525), .in_5 (n_27526), .in_6 (n_27527), .in_7
       (n_27528), .z (arIll[11]));
  fx68k_mux_1529 mux_arIll_1912_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27633));
  fx68k_mux_1529 mux_arIll_1929_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27634));
  fx68k_mux_1529 mux_arIll_1946_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27635));
  fx68k_mux_1529 mux_arIll_1963_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27636));
  fx68k_mux_1529 mux_arIll_1980_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27637));
  fx68k_mux_1529 mux_arIll_1997_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27638));
  fx68k_mux_1529 mux_arIll_2014_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b1), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27639));
  fx68k_mux_1529 mux_arIll_2031_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27640));
  fx68k_bmux_1619 mux_arIll_1909_14(.ctl (opcode[8:6]), .in_0
       (n_27633), .in_1 (n_27634), .in_2 (n_27635), .in_3 (n_27636),
       .in_4 (n_27637), .in_5 (n_27638), .in_6 (n_27639), .in_7
       (n_27640), .z (arIll[12]));
  fx68k_mux_1529 mux_arIll_2054_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b1), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27745));
  fx68k_mux_1529 mux_arIll_2071_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27746));
  fx68k_mux_1529 mux_arIll_2088_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27747));
  fx68k_mux_1529 mux_arIll_2105_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27748));
  fx68k_mux_1529 mux_arIll_2122_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27749));
  fx68k_mux_1529 mux_arIll_2139_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27750));
  fx68k_mux_1529 mux_arIll_2156_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b1), .in_10 (1'b1), .in_11
       (1'b1), .in_12 (1'b1), .z (n_27751));
  fx68k_mux_1529 mux_arIll_2173_19(.ctl ({n_26180, n_26181, n_26182,
       n_26183, n_26184, n_26185, n_26186, n_26187, n_26188, n_26189,
       n_26190, n_26191, n_26192}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b0), .in_8 (1'b0), .in_9 (1'b0), .in_10 (1'b0), .in_11
       (1'b0), .in_12 (1'b1), .z (n_27752));
  fx68k_bmux_1619 mux_arIll_2051_14(.ctl (opcode[8:6]), .in_0
       (n_27745), .in_1 (n_27746), .in_2 (n_27747), .in_3 (n_27748),
       .in_4 (n_27749), .in_5 (n_27750), .in_6 (n_27751), .in_7
       (n_27752), .z (arIll[13]));
  CDN_dc logicX_inst(.cf (1'b0), .dcf (1'b1), .z (_X_));
  not g5 (n_101, opcode[11]);
  and g6 (n_27785, n_101, opcode[7]);
  and g7 (n_25122, n_27785, opcode[6]);
  and g1 (n_27768, arIll[0], lineBmap[0]);
  and g38 (n_27769, arIll[1], lineBmap[1]);
  and g39 (n_27770, arIll[2], lineBmap[2]);
  and g40 (n_27771, arIll[3], lineBmap[3]);
  and g41 (n_27772, arIll[4], lineBmap[4]);
  and g42 (n_27773, arIll[5], lineBmap[5]);
  and g44 (n_27775, opcode[8], lineBmap[7]);
  and g45 (n_27776, arIll[8], lineBmap[8]);
  and g46 (n_27777, arIll[9], lineBmap[9]);
  and g48 (n_27779, arIll[11], lineBmap[11]);
  and g49 (n_27780, arIll[12], lineBmap[12]);
  and g50 (n_27781, arIll[13], lineBmap[13]);
  and g51 (n_27782, arIll[14], lineBmap[14]);
  nand g118 (n_27848, n_10, n_73, n_48, opcode[9]);
  nor g8 (n_23477, n_27848, opcode[10]);
  not g122 (n_73, opcode[7]);
  nand g123 (n_27853, n_73, n_10, n_27852);
  not g124 (n_23491, n_27853);
  nand g130 (n_27859, opcode[6], n_73, n_48, opcode[9]);
  nor g132 (n_23501, n_27859, opcode[10]);
  nand g136 (n_27864, n_73, opcode[6], n_27852);
  not g137 (n_23511, n_27864);
  nand g143 (n_27870, n_10, opcode[7], n_48, opcode[9]);
  nor g145 (n_23521, n_27870, opcode[10]);
  nand g153 (n_27878, opcode[10], opcode[11]);
  nor g9 (n_24491, n_27878, n_27879);
  nor g155 (n_27880, opcode[11], opcode[10], opcode[9]);
  nand g156 (n_27882, n_27880, opcode[8]);
  not g157 (n_25804, n_27882);
  not g158 (n_10, opcode[6]);
  not g159 (n_48, opcode[8]);
  nor g161 (n_27852, opcode[11], opcode[10], opcode[8]);
  not g162 (n_33, opcode[9]);
  nand g163 (n_27879, opcode[7], n_48, n_33);
  or g164 (n_27883, n_25512, n_25513);
  or g165 (n_26715, n_25514, n_25515, n_25516, n_27883);
  nor g169 (n_23665, n_8, n_15);
  nand g170 (n_8, n_73, n_7);
  nor g172 (n_7, opcode[8], n_101);
  nand g175 (n_15, n_10, n_14);
  nor g177 (n_14, opcode[10], opcode[9]);
  nor g11 (n_23666, n_8, n_17);
  nand g12 (n_17, n_14, opcode[6]);
  nor g13 (n_23667, n_17, n_19);
  nand g14 (n_19, n_7, opcode[7]);
  nor g15 (n_23668, n_19, n_15);
  nor g16 (n_23669, n_8, n_24);
  nand g17 (n_24, n_10, n_23);
  nor g18 (n_23, n_22, opcode[9]);
  not g19 (n_22, opcode[10]);
  nor g20 (n_23670, n_8, n_26);
  nand g21 (n_26, n_23, opcode[6]);
  nor g22 (n_23671, n_19, n_24);
  nand g23 (n_26440, n_30, n_32);
  nand g24 (n_30, opcode[7], n_29);
  nor g25 (n_29, n_10, n_22);
  nor g26 (n_32, opcode[8], n_31);
  nand g27 (n_31, n_33, opcode[11]);
  nor g211 (n_23682, n_41, n_83, n_125, n_167);
  nor g269 (n_23701, n_23697, n_23698, n_23699, n_23700);
  nor g273 (n_24058, n_27978, n_27981);
  nand g274 (n_27978, n_27977, n_79);
  not g275 (n_27977, movEa[2]);
  not g276 (n_79, movEa[3]);
  nand g277 (n_27981, n_88, n_87);
  not g278 (n_88, movEa[1]);
  not g279 (n_87, movEa[0]);
  nor g280 (n_24059, n_27978, n_27982);
  nand g281 (n_27982, movEa[1], n_87);
  nor g282 (n_24060, n_27978, n_27983);
  nand g283 (n_27983, movEa[1], movEa[0]);
  nor g284 (n_24061, n_27981, n_27984);
  nand g285 (n_27984, movEa[2], n_79);
  nor g286 (n_24062, n_27984, n_27985);
  nand g287 (n_27985, n_88, movEa[0]);
  nor g288 (n_24063, n_27984, n_27982);
  nor g289 (n_24064, n_27984, n_27983);
  nor g290 (n_24065, n_27981, n_27986);
  nand g291 (n_27986, n_27977, movEa[3]);
  nor g300 (n_24352, n_27991, n_27994);
  nand g301 (n_27991, n_87, n_88);
  nand g304 (n_27994, n_79, n_27977);
  nor g307 (n_24353, n_27994, n_27995);
  nand g308 (n_27995, movEa[0], n_88);
  nor g309 (n_24354, n_27994, n_27996);
  nand g310 (n_27996, n_87, movEa[1]);
  nor g311 (n_24355, n_27994, n_27997);
  nand g312 (n_27997, movEa[0], movEa[1]);
  nor g313 (n_24356, n_27991, n_27998);
  nand g314 (n_27998, n_79, movEa[2]);
  nor g315 (n_24357, n_27995, n_27998);
  nor g316 (n_24358, n_27996, n_27998);
  nor g317 (n_24359, n_27997, n_27998);
  nor g318 (n_24360, n_27991, n_27999);
  nand g319 (n_27999, movEa[3], n_27977);
  nor g323 (n_24511, n_153, n_28008);
  nand g324 (n_153, opcode[6], n_152);
  nor g325 (n_152, opcode[10], n_73);
  nand g327 (n_28008, n_33, n_28007);
  nor g329 (n_28007, opcode[11], opcode[8]);
  nor g331 (n_24512, n_28008, n_28011);
  nand g332 (n_28011, opcode[6], n_28010);
  nor g333 (n_28010, n_22, n_73);
  nor g335 (n_24513, n_28011, n_28012);
  nand g336 (n_28012, n_28007, opcode[9]);
  nor g337 (n_24514, n_28015, n_154);
  nand g338 (n_28015, n_10, n_28014);
  nor g340 (n_28014, opcode[10], opcode[7]);
  nand g341 (n_154, n_33, n_28017);
  nor g342 (n_28017, n_101, opcode[8]);
  nor g344 (n_25588, n_154, n_28);
  nand g345 (n_28, n_28014, opcode[6]);
  nor g346 (n_25589, n_154, n_28018);
  nand g347 (n_28018, n_152, n_10);
  nor g348 (n_25590, n_153, n_154);
  nor g349 (n_24515, n_28015, n_28019);
  nand g28 (n_28019, n_28017, opcode[9]);
  nor g29 (n_24516, n_28, n_28019);
  nor g350 (n_24517, n_28018, n_28019);
  nor g31 (n_24518, n_153, n_28019);
  nand g351 (n_24519, n_28022, n_47);
  nand g352 (n_28022, n_28020, n_28021);
  not g353 (n_28020, n_28017);
  nand g354 (n_28021, opcode[6], n_48);
  nor g355 (n_47, n_28025, n_46);
  nor g356 (n_28025, n_28023, n_44);
  nor g357 (n_28023, opcode[9], opcode[10]);
  and g358 (n_28024, opcode[11], n_22);
  and g359 (n_43, n_101, opcode[10]);
  or g360 (n_44, n_28024, n_43);
  nor g361 (n_46, opcode[11], opcode[7]);
  nor g386 (n_24539, n_24536, n_24537, n_24538);
  nand g395 (n_64, n_48, opcode[7], opcode[6]);
  not g400 (n_24619, n_27967);
  not g401 (n_24620, n_27969);
  not g402 (n_24621, n_27964);
  not g403 (n_24622, n_64);
  not g404 (n_41, n_40);
  not g405 (n_83, n_82);
  not g406 (n_167, n_67);
  not g407 (n_125, n_124);
  nor g524 (n_25512, opcode[5], opcode[4]);
  nor g525 (n_25513, opcode[3], n_28159);
  nand g526 (n_28159, n_28158, opcode[4]);
  not g527 (n_28158, opcode[5]);
  nor g528 (n_25514, n_28159, n_28160);
  not g529 (n_28160, opcode[3]);
  nor g530 (n_25515, opcode[3], n_28162);
  nand g531 (n_28162, opcode[5], n_28161);
  not g532 (n_28161, opcode[4]);
  nor g533 (n_25516, n_28162, n_28160);
  nor g534 (n_25517, opcode[3], n_28163);
  nand g535 (n_28163, opcode[5], opcode[4]);
  nor g536 (n_26716, n_28163, n_28160);
  nor g559 (n_25543, n_125, n_167);
  nor g565 (n_26158, n_73, opcode[6]);
  nor g566 (n_26177, n_73, n_10);
  nor g572 (n_26180, n_28226, n_28229);
  nand g573 (n_28226, n_114, n_28225);
  not g574 (n_114, col[1]);
  not g575 (n_28225, col[2]);
  nand g576 (n_28229, n_28227, n_28228);
  not g577 (n_28227, col[0]);
  not g578 (n_28228, col[3]);
  nor g579 (n_26181, n_28226, n_28230);
  nand g580 (n_28230, col[0], n_28228);
  nor g581 (n_26182, n_28229, n_28231);
  nand g582 (n_28231, col[1], n_28225);
  nor g583 (n_26183, n_28231, n_28230);
  nor g584 (n_26184, n_28229, n_28232);
  nand g585 (n_28232, n_114, col[2]);
  nor g586 (n_26185, n_28232, n_28230);
  nor g587 (n_26186, n_28229, n_28233);
  nand g588 (n_28233, col[1], col[2]);
  nor g589 (n_26187, n_28233, n_28230);
  nor g590 (n_26188, n_28226, n_28234);
  nand g591 (n_28234, n_28227, col[3]);
  nor g592 (n_26189, n_28226, n_28235);
  nand g593 (n_28235, col[0], col[3]);
  nor g594 (n_26190, n_28231, n_28234);
  nor g595 (n_26191, n_28231, n_28235);
  nor g596 (n_26192, n_28228, n_28225);
  nor g2457 (n_27105, n_29266, n_29269);
  nand g2458 (n_29266, n_28227, n_114);
  nand g2461 (n_29269, n_28228, n_28225);
  nor g2464 (n_27106, n_29269, n_29270);
  nand g2465 (n_29270, col[0], n_114);
  nor g2466 (n_27107, n_29269, n_29271);
  nand g2467 (n_29271, n_28227, col[1]);
  nor g2468 (n_27108, n_29269, n_29272);
  nand g2469 (n_29272, col[0], col[1]);
  nor g2470 (n_27109, n_29266, n_29273);
  nand g2471 (n_29273, n_28228, col[2]);
  nor g2472 (n_27110, n_29270, n_29273);
  nor g2473 (n_27111, n_29271, n_29273);
  nor g2474 (n_27112, n_29272, n_29273);
  nor g2475 (n_27113, n_29266, n_29274);
  nand g2476 (n_29274, col[3], n_28225);
  nor g2477 (n_27114, n_28228, n_29276);
  nor g2478 (n_29276, col[0], n_29275);
  nand g2479 (n_29275, n_28225, n_114);
  nand g3829 (n_124, opcode[8], opcode[7], opcode[6]);
  nand g3830 (n_40, opcode[8], n_73, n_10);
  nand g3831 (n_82, opcode[8], n_73, opcode[6]);
  nand g3832 (n_67, opcode[8], opcode[7], n_10);
  nand g3833 (n_27963, n_101, n_22);
  nand g3834 (n_27964, n_48, opcode[7], n_10);
  nand g3835 (n_81, n_101, opcode[10]);
  nand g3836 (n_27967, n_48, n_73, n_10);
  nand g3837 (n_27969, n_48, n_73, opcode[6]);
  nor g3838 (n_23697, n_27963, n_27964);
  nor g3839 (n_23698, n_81, n_27967);
  nor g3840 (n_23699, n_81, n_27969);
  nor g3841 (n_23700, n_81, n_27964);
  nor g3842 (n_24536, opcode[11], n_27967);
  nor g3843 (n_24537, opcode[11], n_27969);
  nor g3844 (n_24538, opcode[11], n_27964);
endmodule

module fx68k_equal_unsigned_1672(A, B, Z);
  input [15:0] A;
  input [6:0] B;
  output Z;
  wire [15:0] A;
  wire [6:0] B;
  wire Z;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32;
  wire n_33, n_34, n_35, n_36, n_37;
  xnor g1 (n_26, A[0], B[0]);
  xnor g2 (n_27, A[1], B[1]);
  xnor g3 (n_28, A[2], B[2]);
  xnor g4 (n_29, A[3], B[3]);
  xnor g5 (n_30, A[4], B[4]);
  xnor g6 (n_31, A[5], B[5]);
  xnor g7 (n_32, A[6], B[6]);
  nor g8 (n_33, A[15], A[14], A[13], A[12]);
  nor g9 (n_34, A[11], A[10], A[9], A[8]);
  not g10 (n_25, A[7]);
  nand g11 (n_35, n_25, n_26, n_27, n_28);
  nand g12 (n_36, n_29, n_30, n_31, n_32);
  nand g13 (n_37, n_33, n_34);
  nor g14 (Z, n_35, n_36, n_37);
endmodule

module fx68k_equal_unsigned_1674(A, B, Z);
  input [15:0] A;
  input [14:0] B;
  output Z;
  wire [15:0] A;
  wire [14:0] B;
  wire Z;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_52;
  xnor g1 (n_34, A[0], B[0]);
  xnor g2 (n_35, A[1], B[1]);
  xnor g3 (n_36, A[2], B[2]);
  xnor g4 (n_37, A[3], B[3]);
  xnor g5 (n_38, A[4], B[4]);
  xnor g6 (n_39, A[5], B[5]);
  xnor g7 (n_40, A[6], B[6]);
  xnor g8 (n_41, A[7], B[7]);
  xnor g9 (n_42, A[8], B[8]);
  xnor g10 (n_43, A[9], B[9]);
  xnor g11 (n_44, A[10], B[10]);
  xnor g12 (n_45, A[11], B[11]);
  xnor g13 (n_46, A[12], B[12]);
  xnor g14 (n_47, A[13], B[13]);
  xnor g15 (n_48, A[14], B[14]);
  not g16 (n_33, A[15]);
  nand g17 (n_49, n_33, n_34, n_35, n_36);
  nand g18 (n_50, n_37, n_38, n_39, n_40);
  nand g19 (n_51, n_41, n_42, n_43, n_44);
  nand g20 (n_52, n_45, n_46, n_47, n_48);
  nor g21 (Z, n_49, n_50, n_51, n_52);
endmodule

module fx68k_case_box_989(in_0, out_0);
  input [2:0] in_0;
  output [5:0] out_0;
  wire [2:0] in_0;
  wire [5:0] out_0;
  wire n_5, n_6, n_8, n_10, n_12, n_16, n_40, n_41;
  nor g1 (out_0[5], in_0[2], n_6);
  nand g2 (n_6, n_40, n_5);
  not g3 (n_40, in_0[1]);
  not g4 (n_5, in_0[0]);
  nor g5 (out_0[4], in_0[2], n_8);
  nand g6 (n_8, n_40, in_0[0]);
  nor g7 (out_0[3], in_0[2], n_10);
  nand g8 (n_10, in_0[1], n_5);
  nor g9 (out_0[2], in_0[2], n_12);
  nand g10 (n_12, in_0[1], in_0[0]);
  nor g11 (out_0[1], n_6, n_41);
  not g12 (n_41, in_0[2]);
  nor g13 (out_0[0], n_16, n_41);
  not g14 (n_16, n_6);
endmodule

module fx68k_mux_1665(ctl, in_0, in_1, in_2, in_3, in_4, in_5, z);
  input [5:0] ctl;
  input [3:0] in_0, in_1, in_2, in_3, in_4, in_5;
  output [3:0] z;
  wire [5:0] ctl;
  wire [3:0] in_0, in_1, in_2, in_3, in_4, in_5;
  wire [3:0] z;
  CDN_mux6 g1(.sel0 (ctl[5]), .data0 (in_0[3]), .sel1 (ctl[4]), .data1
       (in_1[3]), .sel2 (ctl[3]), .data2 (in_2[3]), .sel3 (ctl[2]),
       .data3 (in_3[3]), .sel4 (ctl[1]), .data4 (in_4[3]), .sel5
       (ctl[0]), .data5 (in_5[3]), .z (z[3]));
  CDN_mux6 g5(.sel0 (ctl[5]), .data0 (in_0[2]), .sel1 (ctl[4]), .data1
       (in_1[2]), .sel2 (ctl[3]), .data2 (in_2[2]), .sel3 (ctl[2]),
       .data3 (in_3[2]), .sel4 (ctl[1]), .data4 (in_4[2]), .sel5
       (ctl[0]), .data5 (in_5[2]), .z (z[2]));
  CDN_mux6 g6(.sel0 (ctl[5]), .data0 (in_0[1]), .sel1 (ctl[4]), .data1
       (in_1[1]), .sel2 (ctl[3]), .data2 (in_2[1]), .sel3 (ctl[2]),
       .data3 (in_3[1]), .sel4 (ctl[1]), .data4 (in_4[1]), .sel5
       (ctl[0]), .data5 (in_5[1]), .z (z[1]));
  CDN_mux6 g7(.sel0 (ctl[5]), .data0 (in_0[0]), .sel1 (ctl[4]), .data1
       (in_1[0]), .sel2 (ctl[3]), .data2 (in_2[0]), .sel3 (ctl[2]),
       .data3 (in_3[0]), .sel4 (ctl[1]), .data4 (in_4[0]), .sel5
       (ctl[0]), .data5 (in_5[0]), .z (z[0]));
endmodule

module fx68k_mux_1668(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input [3:0] in_0, in_1;
  output [3:0] z;
  wire [1:0] ctl;
  wire [3:0] in_0, in_1;
  wire [3:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[3]), .sel1 (ctl[0]), .data1
       (in_1[3]), .z (z[3]));
  CDN_mux2 g5(.sel0 (ctl[1]), .data0 (in_0[2]), .sel1 (ctl[0]), .data1
       (in_1[2]), .z (z[2]));
  CDN_mux2 g6(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g7(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_uaddrDecode(opcode, a1, a2, a3, isPriv, isIllegal,
     isLineA, isLineF, lineBmap);
  input [15:0] opcode;
  output [9:0] a1, a2, a3;
  output isPriv, isIllegal, isLineA, isLineF;
  output [15:0] lineBmap;
  wire [15:0] opcode;
  wire [9:0] a1, a2, a3;
  wire isPriv, isIllegal, isLineA, isLineF;
  wire [15:0] lineBmap;
  wire [3:0] movEa;
  wire [3:0] eaCol;
  wire [3:0] eaDecode;
  wire \eaDecode[0]_275 , \eaDecode[1]_276 , \eaDecode[2]_277 ,
       \eaDecode[3]_278 , n_17, n_18, n_19, n_20;
  wire n_23, n_28, n_33, n_36, n_38, n_39, n_40, n_43;
  wire n_48, n_53, n_136, n_137, n_138, n_139, n_140, n_157;
  wire n_158, n_159, n_160, n_161, n_174, n_175, n_176, n_177;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_269, n_270, n_271, n_272, n_273, n_274, n_279, n_280;
  wire n_284, n_285, n_286, n_288, n_289, n_290, n_292, n_293;
  assign lineBmap[10] = isLineA;
  assign lineBmap[15] = isLineF;
  fx68k_onehotEncoder4 irLineDecod(opcode[15:12], {isLineF,
       lineBmap[14:11], isLineA, lineBmap[9:0]});
  fx68k_pla_lined pla_lined(.movEa (movEa), .col (eaCol), .opcode
       (opcode), .lineBmap ({isLineF, lineBmap[14:11], isLineA,
       lineBmap[9:0]}), .palIll (isIllegal), .plaA1 (a1), .plaA2 (a2),
       .plaA3 (a3));
  fx68k_equal_unsigned_1672 eq_1836_41(.A ({opcode[15:12], 1'b0,
       opcode[10], 1'b0, opcode[8:0]}), .B (7'b1111100), .Z (n_160));
  fx68k_equal_unsigned_1674 eq_1841_29(.A ({opcode[15:6], 6'b000000}),
       .B (15'b100011011000000), .Z (n_136));
  fx68k_equal_unsigned_1674 eq_1844_34(.A ({opcode[15:4], 4'b0000}), .B
       (15'b100111001100000), .Z (n_137));
  fx68k_equal_unsigned_1674 eq_1847_21(.A (opcode), .B
       (15'b100111001110000), .Z (n_174));
  fx68k_equal_unsigned_1674 eq_1848_15(.A (opcode), .B
       (15'b100111001110011), .Z (n_175));
  fx68k_equal_unsigned_1674 eq_1849_15(.A (opcode), .B
       (15'b100111001110010), .Z (n_177));
  fx68k_bmux_1503 mux_isPriv_1848_27(.ctl (n_138), .in_0 (1'b0), .in_1
       (1'b1), .z (n_139));
  fx68k_bmux_1503 mux_isPriv_1844_34(.ctl (n_137), .in_0 (n_139), .in_1
       (1'b1), .z (n_140));
  fx68k_bmux_1503 mux_isPriv_1841_29(.ctl (n_136), .in_0 (n_140), .in_1
       (1'b1), .z (n_161));
  fx68k_mux_1527 mux_isPriv_1833_16(.ctl ({n_157, n_158, n_159}), .in_0
       (n_160), .in_1 (n_161), .in_2 (1'b0), .z (isPriv));
  fx68k_case_box_989 ctl_eaBits_1806_9(.in_0 (opcode[2:0]), .out_0
       ({n_258, n_259, n_260, n_261, n_262, n_263}));
  fx68k_mux_1665 \eaDecode_1797_17:mux_eaDecode_1806_9 (.ctl ({n_258,
       n_259, n_260, n_261, n_262, n_263}), .in_0 (4'b0111), .in_1
       (4'b1000), .in_2 (4'b1001), .in_3 (4'b1010), .in_4 (4'b1011),
       .in_5 (4'b1100), .z (eaDecode));
  fx68k_mux_1668 \eaDecode_1797_17:mux_eaDecode_1804_15 (.ctl ({n_264,
       n_265}), .in_0 (eaDecode), .in_1 ({1'b0, opcode[5:3]}), .z
       (eaCol));
  fx68k_case_box_989 ctl_eaBits_1806_10(.in_0 (opcode[11:9]), .out_0
       ({n_269, n_270, n_271, n_272, n_273, n_274}));
  fx68k_mux_1665 \eaDecode_1798_17:mux_eaDecode_1806_9 (.ctl ({n_269,
       n_270, n_271, n_272, n_273, n_274}), .in_0 (4'b0111), .in_1
       (4'b1000), .in_2 (4'b1001), .in_3 (4'b1010), .in_4 (4'b1011),
       .in_5 (4'b1100), .z ({\eaDecode[3]_278 , \eaDecode[2]_277 ,
       \eaDecode[1]_276 , \eaDecode[0]_275 }));
  fx68k_mux_1668 \eaDecode_1798_17:mux_eaDecode_1804_15 (.ctl ({n_279,
       n_280}), .in_0 ({\eaDecode[3]_278 , \eaDecode[2]_277 ,
       \eaDecode[1]_276 , \eaDecode[0]_275 }), .in_1 ({1'b0,
       opcode[8:6]}), .z (movEa));
  or g54 (n_176, n_174, n_175);
  or g55 (n_138, n_176, n_177);
  not g33 (n_284, isLineF);
  not g34 (n_285, lineBmap[14]);
  not g35 (n_286, lineBmap[13]);
  not g36 (n_18, lineBmap[12]);
  not g37 (n_23, lineBmap[11]);
  not g38 (n_28, isLineA);
  not g39 (n_33, lineBmap[9]);
  not g40 (n_38, lineBmap[8]);
  not g41 (n_43, lineBmap[7]);
  not g42 (n_48, lineBmap[6]);
  not g43 (n_53, lineBmap[5]);
  not g45 (n_288, lineBmap[3]);
  not g46 (n_289, lineBmap[2]);
  not g47 (n_290, lineBmap[1]);
  nand g1 (n_17, n_284, n_285, n_286, n_18);
  nand g2 (n_293, n_23, n_28, n_33, n_38);
  nand g3 (n_19, n_43, n_48, n_53, n_292);
  nand g4 (n_20, n_288, n_289, n_290, lineBmap[0]);
  nor g5 (n_157, n_17, n_293, n_19, n_20);
  nand g8 (n_39, n_43, n_48, n_53, lineBmap[4]);
  nand g9 (n_40, n_288, n_289, n_290, n_36);
  nor g10 (n_158, n_17, n_293, n_39, n_40);
  nor g11 (n_159, n_158, n_157);
  not g12 (n_292, lineBmap[4]);
  not g13 (n_36, lineBmap[0]);
  not g56 (n_264, n_265);
  nand g58 (n_265, opcode[5], opcode[4], opcode[3]);
  not g60 (n_279, n_280);
  nand g62 (n_280, opcode[8], opcode[7], opcode[6]);
endmodule

module fx68k_case_box_1015(in_0, out_0);
  input [1:0] in_0;
  output [2:0] out_0;
  wire [1:0] in_0;
  wire [2:0] out_0;
  wire n_4;
  assign out_0[0] = in_0[0];
  nor g1 (out_0[2], in_0[0], in_0[1]);
  nor g2 (out_0[1], in_0[0], n_4);
  not g3 (n_4, in_0[1]);
endmodule

module fx68k_mux_1694(ctl, in_0, in_1, in_2, z);
  input [2:0] ctl;
  input [1:0] in_0, in_1, in_2;
  output [1:0] z;
  wire [2:0] ctl;
  wire [1:0] in_0, in_1, in_2;
  wire [1:0] z;
  CDN_mux3 g1(.sel0 (ctl[2]), .data0 (in_0[1]), .sel1 (ctl[1]), .data1
       (in_1[1]), .sel2 (ctl[0]), .data2 (in_2[1]), .z (z[1]));
  CDN_mux3 g3(.sel0 (ctl[2]), .data0 (in_0[0]), .sel1 (ctl[1]), .data1
       (in_1[0]), .sel2 (ctl[0]), .data2 (in_2[0]), .z (z[0]));
endmodule

module fx68k_case_box_1016(in_0, out_0);
  input [1:0] in_0;
  output [2:0] out_0;
  wire [1:0] in_0;
  wire [2:0] out_0;
  wire n_23;
  not g1 (out_0[2], in_0[0]);
  nor g2 (out_0[1], out_0[2], in_0[1]);
  nor g3 (out_0[0], out_0[2], n_23);
  not g4 (n_23, in_0[1]);
endmodule

module fx68k_case_box_1019(in_0, out_0);
  input [3:0] in_0;
  output [3:0] out_0;
  wire [3:0] in_0;
  wire [3:0] out_0;
  wire n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13;
  wire n_14, n_16, n_17, n_18, n_19, n_22, n_45, n_74;
  assign out_0[0] = in_0[3];
  not g33 (n_45, in_0[3]);
  nor g1 (out_0[3], in_0[3], n_14);
  nand g3 (n_14, n_11, n_13);
  nand g4 (n_11, in_0[2], n_10);
  not g5 (n_7, in_0[1]);
  not g6 (n_6, in_0[0]);
  and g7 (n_8, in_0[1], n_6);
  and g8 (n_9, n_7, in_0[0]);
  or g9 (n_10, n_8, n_9);
  nand g10 (n_13, in_0[1], n_12);
  not g11 (n_12, in_0[2]);
  nor g12 (out_0[2], n_18, n_74);
  and g13 (n_16, in_0[1], in_0[2]);
  and g14 (n_17, n_7, n_12);
  or g15 (n_18, n_16, n_17);
  nand g16 (n_74, n_45, n_19);
  nand g17 (n_19, n_6, in_0[2]);
  nor g18 (out_0[1], n_19, n_22);
  nand g19 (n_22, in_0[1], n_45);
endmodule

module fx68k_mux_1696(ctl, in_0, in_1, in_2, in_3, z);
  input [3:0] ctl;
  input [1:0] in_0, in_1, in_2, in_3;
  output [1:0] z;
  wire [3:0] ctl;
  wire [1:0] in_0, in_1, in_2, in_3;
  wire [1:0] z;
  CDN_mux4 g1(.sel0 (ctl[3]), .data0 (in_0[1]), .sel1 (ctl[2]), .data1
       (in_1[1]), .sel2 (ctl[1]), .data2 (in_2[1]), .sel3 (ctl[0]),
       .data3 (in_3[1]), .z (z[1]));
  CDN_mux4 g3(.sel0 (ctl[3]), .data0 (in_0[0]), .sel1 (ctl[2]), .data1
       (in_1[0]), .sel2 (ctl[1]), .data2 (in_2[0]), .sel3 (ctl[0]),
       .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_bmux_1705(ctl, in_0, in_1, in_2, in_3, z);
  input [1:0] ctl;
  input in_0, in_1, in_2, in_3;
  output z;
  wire [1:0] ctl;
  wire in_0, in_1, in_2, in_3;
  wire z;
  CDN_bmux4 g1(.sel0 (ctl[0]), .data0 (in_0), .data1 (in_1), .sel1
       (ctl[1]), .data2 (in_2), .data3 (in_3), .z (z));
endmodule

module fx68k_bmux_1706(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16,
     in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25,
     in_26, in_27, in_28, in_29, in_30, z);
  input [4:0] ctl;
  input [1:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17,
       in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26,
       in_27, in_28, in_29, in_30;
  output [1:0] z;
  wire [4:0] ctl;
  wire [1:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17,
       in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26,
       in_27, in_28, in_29, in_30;
  wire [1:0] z;
  CDN_bmux31 g1(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .sel3 (ctl[3]), .data8 (in_8[1]), .data9
       (in_9[1]), .data10 (in_10[1]), .data11 (in_11[1]), .data12
       (in_12[1]), .data13 (in_13[1]), .data14 (in_14[1]), .data15
       (in_15[1]), .sel4 (ctl[4]), .data16 (in_16[1]), .data17
       (in_17[1]), .data18 (in_18[1]), .data19 (in_19[1]), .data20
       (in_20[1]), .data21 (in_21[1]), .data22 (in_22[1]), .data23
       (in_23[1]), .data24 (in_24[1]), .data25 (in_25[1]), .data26
       (in_26[1]), .data27 (in_27[1]), .data28 (in_28[1]), .data29
       (in_29[1]), .data30 (in_30[1]), .z (z[1]));
  CDN_bmux31 g2(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .sel3 (ctl[3]), .data8 (in_8[0]), .data9
       (in_9[0]), .data10 (in_10[0]), .data11 (in_11[0]), .data12
       (in_12[0]), .data13 (in_13[0]), .data14 (in_14[0]), .data15
       (in_15[0]), .sel4 (ctl[4]), .data16 (in_16[0]), .data17
       (in_17[0]), .data18 (in_18[0]), .data19 (in_19[0]), .data20
       (in_20[0]), .data21 (in_21[0]), .data22 (in_22[0]), .data23
       (in_23[0]), .data24 (in_24[0]), .data25 (in_25[0]), .data26
       (in_26[0]), .data27 (in_27[0]), .data28 (in_28[0]), .data29
       (in_29[0]), .data30 (in_30[0]), .z (z[0]));
endmodule

module fx68k_mux_1707(ctl, in_0, in_1, in_2, in_3, in_4, in_5, z);
  input [5:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5;
  output z;
  wire [5:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5;
  wire z;
  CDN_mux6 g1(.sel0 (ctl[5]), .data0 (in_0), .sel1 (ctl[4]), .data1
       (in_1), .sel2 (ctl[3]), .data2 (in_2), .sel3 (ctl[2]), .data3
       (in_3), .sel4 (ctl[1]), .data4 (in_4), .sel5 (ctl[0]), .data5
       (in_5), .z (z));
endmodule

module fx68k_bmux_1709(ctl, in_0, in_1, in_2, in_3, z);
  input [1:0] ctl;
  input [9:0] in_0, in_1, in_2, in_3;
  output [9:0] z;
  wire [1:0] ctl;
  wire [9:0] in_0, in_1, in_2, in_3;
  wire [9:0] z;
  CDN_bmux4 g1(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .z (z[9]));
  CDN_bmux4 g2(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .z (z[8]));
  CDN_bmux4 g3(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .z (z[7]));
  CDN_bmux4 g4(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .z (z[6]));
  CDN_bmux4 g5(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .z (z[5]));
  CDN_bmux4 g6(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .z (z[4]));
  CDN_bmux4 g7(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .z (z[3]));
  CDN_bmux4 g8(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .z (z[2]));
  CDN_bmux4 g9(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .z (z[1]));
  CDN_bmux4 g10(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_mux_1713(ctl, in_0, in_1, in_2, in_3, in_4, z);
  input [4:0] ctl;
  input [3:0] in_0, in_1, in_2, in_3, in_4;
  output [3:0] z;
  wire [4:0] ctl;
  wire [3:0] in_0, in_1, in_2, in_3, in_4;
  wire [3:0] z;
  CDN_mux5 g1(.sel0 (ctl[4]), .data0 (in_0[3]), .sel1 (ctl[3]), .data1
       (in_1[3]), .sel2 (ctl[2]), .data2 (in_2[3]), .sel3 (ctl[1]),
       .data3 (in_3[3]), .sel4 (ctl[0]), .data4 (in_4[3]), .z (z[3]));
  CDN_mux5 g5(.sel0 (ctl[4]), .data0 (in_0[2]), .sel1 (ctl[3]), .data1
       (in_1[2]), .sel2 (ctl[2]), .data2 (in_2[2]), .sel3 (ctl[1]),
       .data3 (in_3[2]), .sel4 (ctl[0]), .data4 (in_4[2]), .z (z[2]));
  CDN_mux5 g6(.sel0 (ctl[4]), .data0 (in_0[1]), .sel1 (ctl[3]), .data1
       (in_1[1]), .sel2 (ctl[2]), .data2 (in_2[1]), .sel3 (ctl[1]),
       .data3 (in_3[1]), .sel4 (ctl[0]), .data4 (in_4[1]), .z (z[1]));
  CDN_mux5 g7(.sel0 (ctl[4]), .data0 (in_0[0]), .sel1 (ctl[3]), .data1
       (in_1[0]), .sel2 (ctl[2]), .data2 (in_2[0]), .sel3 (ctl[1]),
       .data3 (in_3[0]), .sel4 (ctl[0]), .data4 (in_4[0]), .z (z[0]));
endmodule

module fx68k_sequencer(\Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] ,
     \Clks[extReset] , \Clks[clk] , enT3, microLatch, A0Err, BerrA,
     busAddrErr, Spuria, Avia, Tpend, intPend, isIllegal, isPriv,
     excRst, isLineA, isLineF, psw, prenEmpty, au05z, dcr4, ze, i11,
     alue01, Ird, a1, a2, a3, tvn, nma);
  input \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset]
       , \Clks[clk] , enT3, A0Err, BerrA, busAddrErr, Spuria, Avia,
       Tpend, intPend, isIllegal, isPriv, excRst, isLineA, isLineF,
       prenEmpty, au05z, dcr4, ze, i11;
  input [16:0] microLatch;
  input [15:0] psw, Ird;
  input [1:0] alue01;
  input [9:0] a1, a2, a3;
  output [3:0] tvn;
  output [9:0] nma;
  wire \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset] ,
       \Clks[clk] , enT3, A0Err, BerrA, busAddrErr, Spuria, Avia,
       Tpend, intPend, isIllegal, isPriv, excRst, isLineA, isLineF,
       prenEmpty, au05z, dcr4, ze, i11;
  wire [16:0] microLatch;
  wire [15:0] psw, Ird;
  wire [1:0] alue01;
  wire [9:0] a1, a2, a3;
  wire [3:0] tvn;
  wire [9:0] nma;
  wire [1:0] c0c1;
  wire [9:0] grp1Nma;
  wire [9:0] uNma;
  wire A0Sel, UNCONNECTED425, _X_, a0Rst, ccTest, grp0LatchEn,
       grp1LatchEn, inGrp0Exc;
  wire n_4, n_8, n_9, n_20, n_21, n_22, n_23, n_24;
  wire n_32, n_33, n_34, n_203, n_204, n_206, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_222, n_223, n_224, n_226, n_227, n_229, n_230, n_231;
  wire n_232, n_233, n_236, n_237, n_238, n_243, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_269, n_270, n_271, n_272, n_273, n_284, n_287;
  wire n_290, n_293, n_296, n_299, n_302, n_305, n_308, n_311;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_358, n_359, n_362, n_363, n_369, n_370;
  wire n_374, n_376, n_378, n_379, n_380, n_383, n_385, n_386;
  wire n_389, n_393, n_394, n_404, n_405, n_446, n_450, n_451;
  wire n_452, n_453, n_454, n_455, rAutovec, rExcAdrErr, rExcBusErr,
       rExcRst;
  wire rIllegal, rInterrupt, rLineA, rLineF, rPriv, rSpurious, rTrace;
  fx68k_bmux_1503 mux_a0Rst_2142_7(.ctl (\Clks[extReset] ), .in_0
       (1'b0), .in_1 (1'b1), .z (UNCONNECTED425));
  fx68k_bmux_1503 mux_nma_1947_13(.ctl (inGrp0Exc), .in_0 (1'b1), .in_1
       (1'b0), .z (n_206));
  fx68k_bmux_1520 mux_nma_1945_8(.ctl (a0Rst), .in_0 ({n_206, 1'b1}),
       .in_1 (2'b10), .z ({n_325, n_324}));
  fx68k_bmux_1503 mux_1984_19(.ctl (au05z), .in_0 (1'b1), .in_1 (1'b0),
       .z (n_255));
  fx68k_bmux_1520 mux_1985_19(.ctl (au05z), .in_0 (2'b11), .in_1
       (2'b00), .z ({n_256, n_243}));
  fx68k_case_box_1015 ctl_nz1_1993_10(.in_0 (psw[3:2]), .out_0 ({n_209,
       n_210, n_211}));
  fx68k_mux_1694 mux_c0c1_1993_10(.ctl ({n_209, n_210, n_211}), .in_0
       (2'b10), .in_1 (2'b01), .in_2 (2'b11), .z ({n_257, n_246}));
  fx68k_case_box_1016 ctl_ms0_2006_9(.in_0 ({Ird[8], alue01[0]}),
       .out_0 ({n_212, n_213, n_214}));
  fx68k_mux_1694 mux_c0c1_2006_9(.ctl ({n_212, n_213, n_214}), .in_0
       (2'b11), .in_1 (2'b01), .in_2 (2'b10), .z ({n_259, n_247}));
  fx68k_case_box_1019 ctl_m01_2013_9(.in_0 ({au05z, Ird[8], alue01}),
       .out_0 ({n_215, n_216, n_217, n_218}));
  fx68k_mux_1696 mux_c0c1_2013_9(.ctl ({n_215, n_216, n_217, n_218}),
       .in_0 (2'b11), .in_1 (2'b01), .in_2 (2'b10), .in_3 (2'b00), .z
       ({n_260, n_248}));
  fx68k_bmux_1590 mux_ccTest_2053_16(.ctl (Ird[11:8]), .in_0 (1'b1),
       .in_1 (1'b0), .in_2 (n_222), .in_3 (n_223), .in_4 (n_224), .in_5
       (psw[0]), .in_6 (n_226), .in_7 (psw[2]), .in_8 (n_227), .in_9
       (psw[1]), .in_10 (n_229), .in_11 (psw[3]), .in_12 (n_230),
       .in_13 (n_231), .in_14 (n_232), .in_15 (n_233), .z (ccTest));
  fx68k_bmux_1503 mux_2021_19(.ctl (ccTest), .in_0 (1'b0), .in_1
       (1'b1), .z (n_261));
  fx68k_bmux_1503 mux_2022_19(.ctl (ccTest), .in_0 (1'b0), .in_1
       (1'b1), .z (n_249));
  fx68k_bmux_1503 mux_2025_18(.ctl (dcr4), .in_0 (1'b1), .in_1 (1'b0),
       .z (n_262));
  fx68k_bmux_1503 mux_2026_18(.ctl (dcr4), .in_0 (1'b1), .in_1 (1'b0),
       .z (n_250));
  fx68k_bmux_1520 mux_2029_18(.ctl (ze), .in_0 (2'b00), .in_1 (2'b11),
       .z ({n_263, n_251}));
  fx68k_bmux_1520 mux_2032_22(.ctl (n_236), .in_0 (2'b11), .in_1
       (2'b00), .z ({n_264, n_252}));
  fx68k_mux_1527 mux_c0c1_2039_10(.ctl ({n_237, n_238, prenEmpty}),
       .in_0 (1'b1), .in_1 (1'b1), .in_2 (1'b0), .z (n_265));
  fx68k_bmux_1705 mux_c0c1_2039_86(.ctl ({Ird[6], prenEmpty}), .in_0
       (1'b0), .in_1 (microLatch[6]), .in_2 (1'b1), .in_3
       (microLatch[6]), .z (n_254));
  fx68k_bmux_1706 mux_c0c1_1981_16(.ctl (microLatch[6:2]), .in_0 ({i11,
       i11}), .in_1 ({n_255, 1'b1}), .in_2 ({1'b0, n_224}), .in_3
       ({psw[2], psw[2]}), .in_4 ({n_257, n_246}), .in_5 ({psw[3],
       1'b1}), .in_6 ({n_258, 1'b1}), .in_7 ({n_259, n_247}), .in_8
       ({n_260, n_248}), .in_9 ({n_261, 1'b1}), .in_10 ({n_263,
       n_251}), .in_11 ({n_264, n_252}), .in_12 ({n_262, 1'b1}), .in_13
       ({n_227, n_227}), .in_14 ({n_265, n_254}), .in_15 ({_X_, _X_}),
       .in_16 ({_X_, _X_}), .in_17 ({n_256, n_243}), .in_18 ({1'b1,
       n_224}), .in_19 ({_X_, _X_}), .in_20 ({_X_, _X_}), .in_21
       ({1'b1, psw[3]}), .in_22 ({_X_, _X_}), .in_23 ({_X_, _X_}),
       .in_24 ({_X_, _X_}), .in_25 ({1'b1, n_249}), .in_26 ({_X_,
       _X_}), .in_27 ({_X_, _X_}), .in_28 ({1'b1, n_250}), .in_29
       ({_X_, _X_}), .in_30 ({n_265, n_254}), .z (c0c1));
  fx68k_mux_1707 mux_grp1Nma_2113_7(.ctl ({rExcRst, n_269, n_270,
       n_271, n_272, n_273}), .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0),
       .in_3 (1'b0), .in_4 (1'b1), .in_5 (1'b0), .z (grp1Nma[2]));
  fx68k_bmux_299 mux_1963_16(.ctl (A0Sel), .in_0 (a1), .in_1
       ({7'b0111000, grp1Nma[2], 2'b00}), .z ({n_311, n_308, n_305,
       n_302, n_299, n_296, n_293, n_290, n_287, n_284}));
  fx68k_bmux_1709 mux_uNma_1961_10(.ctl (microLatch[3:2]), .in_0
       ({microLatch[14:13], microLatch[6:5], microLatch[10:7],
       microLatch[12:11]}), .in_1 ({n_311, n_308, n_305, n_302, n_299,
       n_296, n_293, n_290, n_287, n_284}), .in_2 (a2), .in_3 (a3), .z
       ({n_323, n_322, n_321, n_320, n_319, n_318, n_317, n_316, n_315,
       n_314}));
  fx68k_bmux_299 mux_uNma_1958_7(.ctl (microLatch[1]), .in_0 ({n_323,
       n_322, n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314}),
       .in_1 ({microLatch[14:13], c0c1, microLatch[10:7],
       microLatch[12:11]}), .z (uNma));
  fx68k_bmux_299 mux_nma_1944_7(.ctl (A0Err), .in_0 (uNma), .in_1
       ({8'b00000000, n_325, n_324}), .z (nma));
  fx68k_bmux_1503 mux_2120_10(.ctl (rSpurious), .in_0 (1'b1), .in_1
       (1'b0), .z (n_339));
  fx68k_mux_1713 mux_tvn_2129_11(.ctl ({rIllegal, rPriv, rLineA,
       rLineF, n_330}), .in_0 (4'b0100), .in_1 (4'b1000), .in_2
       (4'b1010), .in_3 (4'b1011), .in_4 (4'b0001), .z ({n_334, n_333,
       n_332, n_331}));
  fx68k_bmux_1504 mux_tvn_2124_12(.ctl (rInterrupt), .in_0 ({n_334,
       n_333, n_332, n_331}), .in_1 (4'b1111), .z ({n_338, n_337,
       n_336, n_335}));
  fx68k_bmux_1504 mux_tvn_2122_12(.ctl (rTrace), .in_0 ({n_338, n_337,
       n_336, n_335}), .in_1 (4'b1001), .z ({n_343, n_342, n_341,
       n_340}));
  fx68k_bmux_1504 mux_tvn_2119_22(.ctl (n_9), .in_0 ({n_343, n_342,
       n_341, n_340}), .in_1 ({3'b110, n_339}), .z ({n_347, n_346,
       n_345, n_344}));
  fx68k_bmux_1504 mux_tvn_2115_23(.ctl (n_8), .in_0 ({n_347, n_346,
       n_345, n_344}), .in_1 ({3'b001, rExcAdrErr}), .z ({n_351, n_350,
       n_349, n_348}));
  fx68k_bmux_1504 mux_tvn_2113_7(.ctl (rExcRst), .in_0 ({n_351, n_350,
       n_349, n_348}), .in_1 (4'b0000), .z (tvn));
  not g1 (n_224, psw[0]);
  not g3 (n_229, psw[3]);
  not g4 (n_226, psw[2]);
  and g5 (n_258, n_229, n_226);
  not g6 (n_227, psw[1]);
  and g9 (n_222, n_224, n_226);
  or g10 (n_223, psw[0], psw[2]);
  and g15 (n_358, psw[3], psw[1]);
  and g18 (n_359, n_229, n_227);
  or g19 (n_230, n_358, n_359);
  and g21 (n_362, psw[3], n_227);
  and g23 (n_363, n_229, psw[1]);
  or g24 (n_231, n_362, n_363);
  and g27 (n_369, n_358, n_226);
  and g31 (n_370, n_359, n_226);
  or g32 (n_232, n_369, n_370);
  or g35 (n_374, psw[2], n_362);
  or g38 (n_233, n_374, n_363);
  or g40 (n_378, microLatch[1], n_376);
  and g41 (grp1LatchEn, microLatch[0], n_378);
  and g43 (grp0LatchEn, microLatch[4], n_379);
  or g44 (n_380, rExcRst, rExcBusErr);
  or g45 (inGrp0Exc, n_380, rExcAdrErr);
  and g46 (n_203, grp0LatchEn, enT3);
  and g47 (n_204, grp1LatchEn, enT3);
  not g48 (n_383, isLineA);
  and g49 (n_385, isIllegal, n_383);
  not g50 (n_386, isLineF);
  and g51 (n_393, n_385, n_386);
  and g53 (n_394, isPriv, n_389);
  or g65 (n_8, rExcBusErr, rExcAdrErr);
  or g66 (n_9, rSpurious, rAutovec);
  not g73 (n_404, \Clks[extReset] );
  CDN_dc logicX_inst(.cf (1'b0), .dcf (1'b1), .z (_X_));
  and g94 (n_405, enT3, n_404);
  not g95 (n_376, microLatch[4]);
  not g96 (n_379, microLatch[1]);
  not g97 (n_389, psw[13]);
  CDN_flop rTrace_reg(.clk (\Clks[clk] ), .d (Tpend), .sena (n_204),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rTrace));
  CDN_flop rInterrupt_reg(.clk (\Clks[clk] ), .d (intPend), .sena
       (n_204), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (rInterrupt));
  CDN_flop rIllegal_reg(.clk (\Clks[clk] ), .d (n_393), .sena (n_204),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rIllegal));
  CDN_flop rPriv_reg(.clk (\Clks[clk] ), .d (n_394), .sena (n_204),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rPriv));
  CDN_flop rLineA_reg(.clk (\Clks[clk] ), .d (isLineA), .sena (n_204),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rLineA));
  CDN_flop rLineF_reg(.clk (\Clks[clk] ), .d (isLineF), .sena (n_204),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rLineF));
  CDN_flop rExcRst_reg(.clk (\Clks[clk] ), .d (excRst), .sena (n_203),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rExcRst));
  CDN_flop rExcAdrErr_reg(.clk (\Clks[clk] ), .d (busAddrErr), .sena
       (n_203), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (rExcAdrErr));
  CDN_flop rExcBusErr_reg(.clk (\Clks[clk] ), .d (BerrA), .sena
       (n_203), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (rExcBusErr));
  CDN_flop rSpurious_reg(.clk (\Clks[clk] ), .d (Spuria), .sena
       (n_203), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (rSpurious));
  CDN_flop rAutovec_reg(.clk (\Clks[clk] ), .d (Avia), .sena (n_203),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rAutovec));
  CDN_flop a0Rst_reg(.clk (\Clks[clk] ), .d (1'b0), .sena (1'b0), .aclr
       (1'b0), .apre (1'b0), .srl (n_446), .srd (\Clks[extReset] ), .q
       (a0Rst));
  or g109 (n_446, n_405, \Clks[extReset] );
  nand g114 (n_450, n_227, n_229);
  not g115 (n_236, n_450);
  or g116 (n_451, rIllegal, rLineF);
  or g117 (n_452, rLineA, rPriv);
  or g118 (A0Sel, rTrace, rInterrupt, n_451, n_452);
  nor g121 (n_237, prenEmpty, Ird[6]);
  nor g2 (n_238, prenEmpty, n_4);
  not g122 (n_4, Ird[6]);
  or g123 (n_20, n_8, rExcRst);
  or g126 (n_23, n_9, n_20);
  not g127 (n_21, rExcRst);
  and g128 (n_269, n_21, n_8);
  not g7 (n_22, n_20);
  and g8 (n_270, n_22, n_9);
  not g129 (n_24, n_23);
  and g130 (n_271, n_24, rTrace);
  nor g132 (n_32, rExcRst, n_8, n_9, rTrace);
  not g133 (n_33, rInterrupt);
  nand g20 (n_34, n_32, n_33);
  not g134 (n_273, n_34);
  nor g139 (n_330, rIllegal, rPriv, rLineA, rLineF);
  and g140 (n_272, n_453, n_454, n_455, rInterrupt);
  not g141 (n_453, rTrace);
  not g142 (n_454, n_9);
  not g143 (n_455, n_20);
endmodule

module fx68k_case_box_1035(in_0, out_0);
  input [15:0] in_0;
  output [16:0] out_0;
  wire [15:0] in_0;
  wire [16:0] out_0;
  wire n_80, n_93, n_139, n_159, n_169, n_198, n_207, n_218;
  wire n_238, n_245, n_257, n_258, n_297, n_302, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_337, n_338;
  wire n_339, n_340, n_341;
  assign out_0[16] = in_0[0];
  nand g19 (n_80, in_0[3], n_321, n_319, n_317);
  nand g24 (n_323, n_93, n_321, n_319, n_317);
  nand g38 (n_159, in_0[7], n_326, n_325, n_322);
  nand g43 (n_328, n_169, n_326, n_325, n_322);
  nand g57 (n_238, in_0[11], n_329, n_207, n_327);
  nand g62 (n_258, n_245, n_329, n_207, n_327);
  nor g65 (out_0[4], n_257, n_258, n_328, n_323);
  nor g70 (out_0[3], n_330, n_258, n_328, n_323);
  nor g75 (out_0[2], n_297, n_258, n_328, n_323);
  nand g76 (n_332, in_0[15], n_302, n_331, n_257);
  nor g80 (out_0[1], n_332, n_258, n_328, n_323);
  nor g81 (n_337, in_0[0], out_0[15], out_0[14], out_0[13]);
  nor g82 (n_338, out_0[12], out_0[11], out_0[10], out_0[9]);
  nor g83 (n_339, out_0[8], out_0[7], out_0[6], out_0[5]);
  nor g84 (n_340, out_0[4], out_0[3], out_0[2], out_0[1]);
  nand g85 (n_341, n_337, n_338, n_339, n_340);
  not g86 (out_0[0], n_341);
  not g87 (n_317, in_0[0]);
  not g88 (n_319, in_0[1]);
  not g89 (n_321, in_0[2]);
  not g90 (n_93, in_0[3]);
  not g91 (n_322, in_0[4]);
  not g92 (n_325, in_0[5]);
  not g93 (n_326, in_0[6]);
  not g94 (n_169, in_0[7]);
  not g95 (n_327, in_0[8]);
  not g96 (n_207, in_0[9]);
  not g97 (n_329, in_0[10]);
  not g98 (n_245, in_0[11]);
  not g99 (n_257, in_0[12]);
  not g100 (n_331, in_0[13]);
  not g101 (n_302, in_0[14]);
  nand g102 (n_318, in_0[1], n_317);
  nand g103 (n_320, in_0[2], n_319, n_317);
  nand g104 (n_324, in_0[5], n_322);
  nand g105 (n_139, in_0[6], n_325, n_322);
  nand g106 (n_198, in_0[9], n_327);
  nand g107 (n_218, in_0[10], n_207, n_327);
  nand g108 (n_330, in_0[13], n_257);
  nand g109 (n_297, in_0[14], n_331, n_257);
  not g110 (out_0[15], n_318);
  not g111 (out_0[14], n_320);
  not g112 (out_0[13], n_80);
  nor g113 (out_0[12], n_322, n_323);
  nor g114 (out_0[11], n_324, n_323);
  nor g115 (out_0[10], n_139, n_323);
  nor g116 (out_0[9], n_159, n_323);
  nor g117 (out_0[8], n_327, n_328, n_323);
  nor g118 (out_0[7], n_198, n_328, n_323);
  nor g119 (out_0[6], n_218, n_328, n_323);
  nor g120 (out_0[5], n_238, n_328, n_323);
endmodule

module fx68k_mux_1721(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16,
     z);
  input [16:0] ctl;
  input [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16;
  output [3:0] z;
  wire [16:0] ctl;
  wire [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16;
  wire [3:0] z;
  CDN_mux17 g1(.sel0 (ctl[16]), .data0 (in_0[3]), .sel1 (ctl[15]),
       .data1 (in_1[3]), .sel2 (ctl[14]), .data2 (in_2[3]), .sel3
       (ctl[13]), .data3 (in_3[3]), .sel4 (ctl[12]), .data4 (in_4[3]),
       .sel5 (ctl[11]), .data5 (in_5[3]), .sel6 (ctl[10]), .data6
       (in_6[3]), .sel7 (ctl[9]), .data7 (in_7[3]), .sel8 (ctl[8]),
       .data8 (in_8[3]), .sel9 (ctl[7]), .data9 (in_9[3]), .sel10
       (ctl[6]), .data10 (in_10[3]), .sel11 (ctl[5]), .data11
       (in_11[3]), .sel12 (ctl[4]), .data12 (in_12[3]), .sel13
       (ctl[3]), .data13 (in_13[3]), .sel14 (ctl[2]), .data14
       (in_14[3]), .sel15 (ctl[1]), .data15 (in_15[3]), .sel16
       (ctl[0]), .data16 (in_16[3]), .z (z[3]));
  CDN_mux17 g5(.sel0 (ctl[16]), .data0 (in_0[2]), .sel1 (ctl[15]),
       .data1 (in_1[2]), .sel2 (ctl[14]), .data2 (in_2[2]), .sel3
       (ctl[13]), .data3 (in_3[2]), .sel4 (ctl[12]), .data4 (in_4[2]),
       .sel5 (ctl[11]), .data5 (in_5[2]), .sel6 (ctl[10]), .data6
       (in_6[2]), .sel7 (ctl[9]), .data7 (in_7[2]), .sel8 (ctl[8]),
       .data8 (in_8[2]), .sel9 (ctl[7]), .data9 (in_9[2]), .sel10
       (ctl[6]), .data10 (in_10[2]), .sel11 (ctl[5]), .data11
       (in_11[2]), .sel12 (ctl[4]), .data12 (in_12[2]), .sel13
       (ctl[3]), .data13 (in_13[2]), .sel14 (ctl[2]), .data14
       (in_14[2]), .sel15 (ctl[1]), .data15 (in_15[2]), .sel16
       (ctl[0]), .data16 (in_16[2]), .z (z[2]));
  CDN_mux17 g6(.sel0 (ctl[16]), .data0 (in_0[1]), .sel1 (ctl[15]),
       .data1 (in_1[1]), .sel2 (ctl[14]), .data2 (in_2[1]), .sel3
       (ctl[13]), .data3 (in_3[1]), .sel4 (ctl[12]), .data4 (in_4[1]),
       .sel5 (ctl[11]), .data5 (in_5[1]), .sel6 (ctl[10]), .data6
       (in_6[1]), .sel7 (ctl[9]), .data7 (in_7[1]), .sel8 (ctl[8]),
       .data8 (in_8[1]), .sel9 (ctl[7]), .data9 (in_9[1]), .sel10
       (ctl[6]), .data10 (in_10[1]), .sel11 (ctl[5]), .data11
       (in_11[1]), .sel12 (ctl[4]), .data12 (in_12[1]), .sel13
       (ctl[3]), .data13 (in_13[1]), .sel14 (ctl[2]), .data14
       (in_14[1]), .sel15 (ctl[1]), .data15 (in_15[1]), .sel16
       (ctl[0]), .data16 (in_16[1]), .z (z[1]));
  CDN_mux17 g7(.sel0 (ctl[16]), .data0 (in_0[0]), .sel1 (ctl[15]),
       .data1 (in_1[0]), .sel2 (ctl[14]), .data2 (in_2[0]), .sel3
       (ctl[13]), .data3 (in_3[0]), .sel4 (ctl[12]), .data4 (in_4[0]),
       .sel5 (ctl[11]), .data5 (in_5[0]), .sel6 (ctl[10]), .data6
       (in_6[0]), .sel7 (ctl[9]), .data7 (in_7[0]), .sel8 (ctl[8]),
       .data8 (in_8[0]), .sel9 (ctl[7]), .data9 (in_9[0]), .sel10
       (ctl[6]), .data10 (in_10[0]), .sel11 (ctl[5]), .data11
       (in_11[0]), .sel12 (ctl[4]), .data12 (in_12[0]), .sel13
       (ctl[3]), .data13 (in_13[0]), .sel14 (ctl[2]), .data14
       (in_14[0]), .sel15 (ctl[1]), .data15 (in_15[0]), .sel16
       (ctl[0]), .data16 (in_16[0]), .z (z[0]));
endmodule

module fx68k_pren(mask, hbit);
  input [15:0] mask;
  output [3:0] hbit;
  wire [15:0] mask;
  wire [3:0] hbit;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101;
  fx68k_case_box_1035 ctl_mask_1903_15(.in_0 (mask), .out_0 ({n_85,
       n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95,
       n_96, n_97, n_98, n_99, n_100, n_101}));
  fx68k_mux_1721 mux_hbit_1903_15(.ctl ({n_85, n_86, n_87, n_88, n_89,
       n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99,
       n_100, n_101}), .in_0 (4'b0000), .in_1 (4'b0001), .in_2
       (4'b0010), .in_3 (4'b0011), .in_4 (4'b0100), .in_5 (4'b0101),
       .in_6 (4'b0110), .in_7 (4'b0111), .in_8 (4'b1000), .in_9
       (4'b1001), .in_10 (4'b1010), .in_11 (4'b1011), .in_12 (4'b1100),
       .in_13 (4'b1101), .in_14 (4'b1110), .in_15 (4'b1111), .in_16
       (4'b0000), .z (hbit));
endmodule

module fx68k_dataIo(\Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] ,
     \Clks[extReset] , \Clks[clk] , enT1, enT2, enT3, enT4,
     \Nanod[abdIsByte] , \Nanod[dblDbh] , \Nanod[dblDbd] ,
     \Nanod[ablAbh] , \Nanod[ablAbd] , \Nanod[extAbh] , \Nanod[extDbh]
     , \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] , \Nanod[au2Pc] ,
     \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd] , \Nanod[alu2Dbd]
     , \Nanod[abd2Alub] , \Nanod[dbd2Alub] , \Nanod[alue2Dbd] ,
     \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] , \Nanod[abd2Dcr] ,
     \Nanod[aluFinish] , \Nanod[aluInit] , \Nanod[aluActrl] ,
     \Nanod[aluDctrl] , \Nanod[aluColumn] , \Nanod[rxlDbl] , \Nanod[rz]
     , \Nanod[abl2ryl] , \Nanod[dbl2ryl] , \Nanod[ryh2abh] ,
     \Nanod[ryh2dbh] , \Nanod[ryl2ab] , \Nanod[ryl2db] ,
     \Nanod[abh2ryh] , \Nanod[dbh2ryh] , \Nanod[abh2rxh] ,
     \Nanod[abl2rxl] , \Nanod[rxl2ab] , \Nanod[rxl2db] ,
     \Nanod[dbh2rxh] , \Nanod[dbl2rxl] , \Nanod[rxh2abh] ,
     \Nanod[rxh2dbh] , \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl]
     , \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
     , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
     \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
     \Nanod[dobCtrl] , \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob]
     , \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
     \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
     \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
     \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] , \Nanod[auCntrl]
     , \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
     \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
     \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
     \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
     \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
     \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
     \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
     \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
     \Nanod[waitBusFinish] , \Nanod[permStart] , \Irdecod[inhibitCcr] ,
     \Irdecod[macroTvn] , \Irdecod[ftuConst] , \Irdecod[ryIsAreg] ,
     \Irdecod[rxIsAreg] , \Irdecod[ry] , \Irdecod[rx] ,
     \Irdecod[isMovep] , \Irdecod[isByte] , \Irdecod[movemPreDecr] ,
     \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] ,
     \Irdecod[rxIsDt] , \Irdecod[toCcr] , \Irdecod[implicitSp] ,
     \Irdecod[isTas] , \Irdecod[isPcRel] , iEdb, aob0, dobIdle,
     dobInput, Irc, dbin, oEdb);
  input \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset]
       , \Clks[clk] , enT1, enT2, enT3, enT4, \Nanod[abdIsByte] ,
       \Nanod[dblDbh] , \Nanod[dblDbd] , \Nanod[ablAbh] ,
       \Nanod[ablAbd] , \Nanod[extAbh] , \Nanod[extDbh] ,
       \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] , \Nanod[au2Pc] ,
       \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd] ,
       \Nanod[alu2Dbd] , \Nanod[abd2Alub] , \Nanod[dbd2Alub] ,
       \Nanod[alue2Dbd] , \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] ,
       \Nanod[abd2Dcr] , \Nanod[aluFinish] , \Nanod[aluInit] ,
       \Nanod[aluActrl] , \Nanod[rxlDbl] , \Nanod[rz] , \Nanod[abl2ryl]
       , \Nanod[dbl2ryl] , \Nanod[ryh2abh] , \Nanod[ryh2dbh] ,
       \Nanod[ryl2ab] , \Nanod[ryl2db] , \Nanod[abh2ryh] ,
       \Nanod[dbh2ryh] , \Nanod[abh2rxh] , \Nanod[abl2rxl] ,
       \Nanod[rxl2ab] , \Nanod[rxl2db] , \Nanod[dbh2rxh] ,
       \Nanod[dbl2rxl] , \Nanod[rxh2abh] , \Nanod[rxh2dbh] ,
       \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl] ,
       \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
       , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
       \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
       \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob] ,
       \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
       \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
       \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
       \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] ,
       \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
       \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
       \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
       \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
       \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
       \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
       \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
       \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
       \Nanod[waitBusFinish] , \Nanod[permStart] , \Irdecod[inhibitCcr]
       , \Irdecod[ryIsAreg] , \Irdecod[rxIsAreg] , \Irdecod[isMovep] ,
       \Irdecod[isByte] , \Irdecod[movemPreDecr] , \Irdecod[rxIsMovem]
       , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] , \Irdecod[rxIsDt] ,
       \Irdecod[toCcr] , \Irdecod[implicitSp] , \Irdecod[isTas] ,
       \Irdecod[isPcRel] , aob0, dobIdle;
  input [1:0] \Nanod[aluDctrl] , \Nanod[dobCtrl] ;
  input [2:0] \Nanod[aluColumn] , \Nanod[auCntrl] , \Irdecod[ry] ,
       \Irdecod[rx] ;
  input [5:0] \Irdecod[macroTvn] ;
  input [15:0] \Irdecod[ftuConst] , iEdb, dobInput;
  output [15:0] Irc, dbin, oEdb;
  wire \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset] ,
       \Clks[clk] , enT1, enT2, enT3, enT4, \Nanod[abdIsByte] ,
       \Nanod[dblDbh] , \Nanod[dblDbd] , \Nanod[ablAbh] ,
       \Nanod[ablAbd] , \Nanod[extAbh] , \Nanod[extDbh] ,
       \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] , \Nanod[au2Pc] ,
       \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd] ,
       \Nanod[alu2Dbd] , \Nanod[abd2Alub] , \Nanod[dbd2Alub] ,
       \Nanod[alue2Dbd] , \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] ,
       \Nanod[abd2Dcr] , \Nanod[aluFinish] , \Nanod[aluInit] ,
       \Nanod[aluActrl] , \Nanod[rxlDbl] , \Nanod[rz] , \Nanod[abl2ryl]
       , \Nanod[dbl2ryl] , \Nanod[ryh2abh] , \Nanod[ryh2dbh] ,
       \Nanod[ryl2ab] , \Nanod[ryl2db] , \Nanod[abh2ryh] ,
       \Nanod[dbh2ryh] , \Nanod[abh2rxh] , \Nanod[abl2rxl] ,
       \Nanod[rxl2ab] , \Nanod[rxl2db] , \Nanod[dbh2rxh] ,
       \Nanod[dbl2rxl] , \Nanod[rxh2abh] , \Nanod[rxh2dbh] ,
       \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl] ,
       \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
       , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
       \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
       \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob] ,
       \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
       \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
       \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
       \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] ,
       \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
       \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
       \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
       \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
       \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
       \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
       \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
       \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
       \Nanod[waitBusFinish] , \Nanod[permStart] , \Irdecod[inhibitCcr]
       , \Irdecod[ryIsAreg] , \Irdecod[rxIsAreg] , \Irdecod[isMovep] ,
       \Irdecod[isByte] , \Irdecod[movemPreDecr] , \Irdecod[rxIsMovem]
       , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] , \Irdecod[rxIsDt] ,
       \Irdecod[toCcr] , \Irdecod[implicitSp] , \Irdecod[isTas] ,
       \Irdecod[isPcRel] , aob0, dobIdle;
  wire [1:0] \Nanod[aluDctrl] , \Nanod[dobCtrl] ;
  wire [2:0] \Nanod[aluColumn] , \Nanod[auCntrl] , \Irdecod[ry] ,
       \Irdecod[rx] ;
  wire [5:0] \Irdecod[macroTvn] ;
  wire [15:0] \Irdecod[ftuConst] , iEdb, dobInput;
  wire [15:0] Irc, dbin, oEdb;
  wire [15:0] dob;
  wire UNCONNECTED426, UNCONNECTED427, byteCycle, byteMux, dbinNoHigh,
       dbinNoLow, isByte_T4, n_4;
  wire n_22, n_27, n_28, n_29, n_46, n_47, n_50, n_51;
  wire n_53, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_77, n_80, n_81, xToDbin, xToIrc;
  fx68k_bmux mux_1761_16(.ctl (\Nanod[noLowByte] ), .in_0
       (dobInput[7:0]), .in_1 (dobInput[15:8]), .z (dob[7:0]));
  fx68k_bmux mux_1762_28(.ctl (n_22), .in_0 (dobInput[15:8]), .in_1
       (dobInput[7:0]), .z (dob[15:8]));
  fx68k_bmux_1503 mux_xToIrc_1722_7(.ctl (enT1), .in_0 (\Nanod[toIrc]
       ), .in_1 (1'b0), .z (UNCONNECTED426));
  fx68k_bmux_1503 mux_xToDbin_1722_7(.ctl (enT1), .in_0 (\Nanod[todbin]
       ), .in_1 (1'b0), .z (UNCONNECTED427));
  fx68k_bmux mux_1740_19(.ctl (byteMux), .in_0 (iEdb[7:0]), .in_1
       (iEdb[15:8]), .z ({n_66, n_65, n_64, n_63, n_62, n_61, n_60,
       n_58}));
  fx68k_bmux mux_1742_29(.ctl (n_46), .in_0 (iEdb[15:8]), .in_1
       (iEdb[7:0]), .z ({n_75, n_74, n_73, n_72, n_71, n_70, n_69,
       n_67}));
  and g1 (n_50, \Nanod[busByte] , isByte_T4);
  not g2 (n_51, aob0);
  and g3 (n_77, n_50, n_51);
  and g4 (n_47, xToIrc, \Clks[enPhi2] );
  and g5 (n_27, xToDbin, \Clks[enPhi2] );
  not g6 (n_29, dbinNoLow);
  not g7 (n_28, dbinNoHigh);
  not g8 (n_53, byteMux);
  and g9 (n_46, n_53, dbinNoLow);
  and g18 (n_81, \Nanod[busByte] , \Irdecod[isByte] );
  not g19 (n_80, dobIdle);
  and g20 (n_4, enT3, n_80);
  or g21 (n_22, byteCycle, \Nanod[noHighByte] );
  and g39 (n_59, n_29, n_27);
  and g40 (n_68, n_28, n_27);
  CDN_flop \Irc_reg[0] (.clk (\Clks[clk] ), .d (iEdb[0]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[0]));
  CDN_flop \Irc_reg[1] (.clk (\Clks[clk] ), .d (iEdb[1]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[1]));
  CDN_flop \Irc_reg[2] (.clk (\Clks[clk] ), .d (iEdb[2]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[2]));
  CDN_flop \Irc_reg[3] (.clk (\Clks[clk] ), .d (iEdb[3]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[3]));
  CDN_flop \Irc_reg[4] (.clk (\Clks[clk] ), .d (iEdb[4]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[4]));
  CDN_flop \Irc_reg[5] (.clk (\Clks[clk] ), .d (iEdb[5]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[5]));
  CDN_flop \Irc_reg[6] (.clk (\Clks[clk] ), .d (iEdb[6]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[6]));
  CDN_flop \Irc_reg[7] (.clk (\Clks[clk] ), .d (iEdb[7]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[7]));
  CDN_flop \Irc_reg[8] (.clk (\Clks[clk] ), .d (iEdb[8]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[8]));
  CDN_flop \Irc_reg[9] (.clk (\Clks[clk] ), .d (iEdb[9]), .sena (n_47),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[9]));
  CDN_flop \Irc_reg[10] (.clk (\Clks[clk] ), .d (iEdb[10]), .sena
       (n_47), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[10]));
  CDN_flop \Irc_reg[11] (.clk (\Clks[clk] ), .d (iEdb[11]), .sena
       (n_47), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[11]));
  CDN_flop \Irc_reg[12] (.clk (\Clks[clk] ), .d (iEdb[12]), .sena
       (n_47), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[12]));
  CDN_flop \Irc_reg[13] (.clk (\Clks[clk] ), .d (iEdb[13]), .sena
       (n_47), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[13]));
  CDN_flop \Irc_reg[14] (.clk (\Clks[clk] ), .d (iEdb[14]), .sena
       (n_47), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[14]));
  CDN_flop \Irc_reg[15] (.clk (\Clks[clk] ), .d (iEdb[15]), .sena
       (n_47), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Irc[15]));
  CDN_flop \dbin_reg[0] (.clk (\Clks[clk] ), .d (n_58), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[0]));
  CDN_flop \dbin_reg[1] (.clk (\Clks[clk] ), .d (n_60), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[1]));
  CDN_flop \dbin_reg[2] (.clk (\Clks[clk] ), .d (n_61), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[2]));
  CDN_flop \dbin_reg[3] (.clk (\Clks[clk] ), .d (n_62), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[3]));
  CDN_flop \dbin_reg[4] (.clk (\Clks[clk] ), .d (n_63), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[4]));
  CDN_flop \dbin_reg[5] (.clk (\Clks[clk] ), .d (n_64), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[5]));
  CDN_flop \dbin_reg[6] (.clk (\Clks[clk] ), .d (n_65), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[6]));
  CDN_flop \dbin_reg[7] (.clk (\Clks[clk] ), .d (n_66), .sena (n_59),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[7]));
  CDN_flop \dbin_reg[8] (.clk (\Clks[clk] ), .d (n_67), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[8]));
  CDN_flop \dbin_reg[9] (.clk (\Clks[clk] ), .d (n_69), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[9]));
  CDN_flop \dbin_reg[10] (.clk (\Clks[clk] ), .d (n_70), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[10]));
  CDN_flop \dbin_reg[11] (.clk (\Clks[clk] ), .d (n_71), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[11]));
  CDN_flop \dbin_reg[12] (.clk (\Clks[clk] ), .d (n_72), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[12]));
  CDN_flop \dbin_reg[13] (.clk (\Clks[clk] ), .d (n_73), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[13]));
  CDN_flop \dbin_reg[14] (.clk (\Clks[clk] ), .d (n_74), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[14]));
  CDN_flop \dbin_reg[15] (.clk (\Clks[clk] ), .d (n_75), .sena (n_68),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dbin[15]));
  CDN_flop xToDbin_reg(.clk (\Clks[clk] ), .d (\Nanod[todbin] ), .sena
       (enT3), .aclr (1'b0), .apre (1'b0), .srl (enT1), .srd (1'b0), .q
       (xToDbin));
  CDN_flop xToIrc_reg(.clk (\Clks[clk] ), .d (\Nanod[toIrc] ), .sena
       (enT3), .aclr (1'b0), .apre (1'b0), .srl (enT1), .srd (1'b0), .q
       (xToIrc));
  CDN_flop dbinNoLow_reg(.clk (\Clks[clk] ), .d (\Nanod[noLowByte] ),
       .sena (enT3), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dbinNoLow));
  CDN_flop dbinNoHigh_reg(.clk (\Clks[clk] ), .d (\Nanod[noHighByte] ),
       .sena (enT3), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dbinNoHigh));
  CDN_flop byteMux_reg(.clk (\Clks[clk] ), .d (n_77), .sena (enT3),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (byteMux));
  CDN_flop isByte_T4_reg(.clk (\Clks[clk] ), .d (\Irdecod[isByte] ),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (isByte_T4));
  CDN_flop \dob_reg[0] (.clk (\Clks[clk] ), .d (dob[0]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[0]));
  CDN_flop \dob_reg[1] (.clk (\Clks[clk] ), .d (dob[1]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[1]));
  CDN_flop \dob_reg[2] (.clk (\Clks[clk] ), .d (dob[2]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[2]));
  CDN_flop \dob_reg[3] (.clk (\Clks[clk] ), .d (dob[3]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[3]));
  CDN_flop \dob_reg[4] (.clk (\Clks[clk] ), .d (dob[4]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[4]));
  CDN_flop \dob_reg[5] (.clk (\Clks[clk] ), .d (dob[5]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[5]));
  CDN_flop \dob_reg[6] (.clk (\Clks[clk] ), .d (dob[6]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[6]));
  CDN_flop \dob_reg[7] (.clk (\Clks[clk] ), .d (dob[7]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[7]));
  CDN_flop \dob_reg[8] (.clk (\Clks[clk] ), .d (dob[8]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[8]));
  CDN_flop \dob_reg[9] (.clk (\Clks[clk] ), .d (dob[9]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[9]));
  CDN_flop \dob_reg[10] (.clk (\Clks[clk] ), .d (dob[10]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[10]));
  CDN_flop \dob_reg[11] (.clk (\Clks[clk] ), .d (dob[11]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[11]));
  CDN_flop \dob_reg[12] (.clk (\Clks[clk] ), .d (dob[12]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[12]));
  CDN_flop \dob_reg[13] (.clk (\Clks[clk] ), .d (dob[13]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[13]));
  CDN_flop \dob_reg[14] (.clk (\Clks[clk] ), .d (dob[14]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[14]));
  CDN_flop \dob_reg[15] (.clk (\Clks[clk] ), .d (dob[15]), .sena (n_4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (oEdb[15]));
  CDN_flop byteCycle_reg(.clk (\Clks[clk] ), .d (n_81), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (byteCycle));
endmodule

module fx68k_case_box_1045(in_0, out_0);
  input [2:0] in_0;
  output [6:0] out_0;
  wire [2:0] in_0;
  wire [6:0] out_0;
  wire n_5, n_6, n_8, n_10, n_13, n_47;
  nor g1 (out_0[6], in_0[0], n_6);
  nand g2 (n_6, n_47, n_5);
  not g3 (n_47, in_0[2]);
  not g4 (n_5, in_0[1]);
  nor g5 (out_0[5], n_6, n_8);
  not g6 (n_8, in_0[0]);
  nor g7 (out_0[4], in_0[0], n_10);
  nand g8 (n_10, n_47, in_0[1]);
  nor g9 (out_0[3], n_10, n_8);
  nor g10 (out_0[2], in_0[0], n_13);
  nand g11 (n_13, in_0[2], n_5);
  nor g12 (out_0[1], n_13, n_8);
  nor g13 (out_0[0], n_47, n_5);
endmodule

module fx68k_mux_1738(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [5:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [5:0] z;
  wire [6:0] ctl;
  wire [5:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [5:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g7(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g8(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g9(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g10(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g11(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_mux_1744(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input [6:0] in_0, in_1;
  output [6:0] z;
  wire [1:0] ctl;
  wire [6:0] in_0, in_1;
  wire [6:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[6]), .sel1 (ctl[0]), .data1
       (in_1[6]), .z (z[6]));
  CDN_mux2 g8(.sel0 (ctl[1]), .data0 (in_0[5]), .sel1 (ctl[0]), .data1
       (in_1[5]), .z (z[5]));
  CDN_mux2 g9(.sel0 (ctl[1]), .data0 (in_0[4]), .sel1 (ctl[0]), .data1
       (in_1[4]), .z (z[4]));
  CDN_mux2 g10(.sel0 (ctl[1]), .data0 (in_0[3]), .sel1 (ctl[0]), .data1
       (in_1[3]), .z (z[3]));
  CDN_mux2 g11(.sel0 (ctl[1]), .data0 (in_0[2]), .sel1 (ctl[0]), .data1
       (in_1[2]), .z (z[2]));
  CDN_mux2 g12(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g13(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_case_box_1049(in_0, out_0);
  input [2:0] in_0;
  output [7:0] out_0;
  wire [2:0] in_0;
  wire [7:0] out_0;
  wire n_5, n_6, n_8, n_10, n_12, n_14, n_54;
  nor g1 (out_0[7], in_0[2], n_6);
  nand g2 (n_6, n_54, n_5);
  not g3 (n_54, in_0[1]);
  not g4 (n_5, in_0[0]);
  nor g5 (out_0[6], in_0[2], n_8);
  nand g6 (n_8, n_54, in_0[0]);
  nor g7 (out_0[5], in_0[2], n_10);
  nand g8 (n_10, in_0[1], n_5);
  nor g9 (out_0[4], in_0[2], n_12);
  nand g10 (n_12, in_0[1], in_0[0]);
  nor g11 (out_0[3], n_6, n_14);
  not g12 (n_14, in_0[2]);
  nor g13 (out_0[2], n_8, n_14);
  nor g14 (out_0[1], n_10, n_14);
  nor g15 (out_0[0], n_12, n_14);
endmodule

module fx68k_mux_1759(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input [5:0] in_0, in_1;
  output [5:0] z;
  wire [1:0] ctl;
  wire [5:0] in_0, in_1;
  wire [5:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[5]), .sel1 (ctl[0]), .data1
       (in_1[5]), .z (z[5]));
  CDN_mux2 g7(.sel0 (ctl[1]), .data0 (in_0[4]), .sel1 (ctl[0]), .data1
       (in_1[4]), .z (z[4]));
  CDN_mux2 g8(.sel0 (ctl[1]), .data0 (in_0[3]), .sel1 (ctl[0]), .data1
       (in_1[3]), .z (z[3]));
  CDN_mux2 g9(.sel0 (ctl[1]), .data0 (in_0[2]), .sel1 (ctl[0]), .data1
       (in_1[2]), .z (z[2]));
  CDN_mux2 g10(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g11(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_bmux_1766(ctl, in_0, in_1, z);
  input ctl;
  input [2:0] in_0, in_1;
  output [2:0] z;
  wire ctl;
  wire [2:0] in_0, in_1;
  wire [2:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_mux_1769(ctl, in_0, in_1, z);
  input [1:0] ctl, in_0, in_1;
  output [1:0] z;
  wire [1:0] ctl, in_0, in_1;
  wire [1:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g3(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_case_box_1064(in_0, out_0);
  input [2:0] in_0;
  output [7:0] out_0;
  wire [2:0] in_0;
  wire [7:0] out_0;
  wire n_25, n_27, n_39, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67;
  nand g1 (n_25, n_60, n_61, n_62);
  nand g2 (n_27, n_60, n_61, in_0[0]);
  nand g3 (n_63, n_60, in_0[1], n_62);
  nand g4 (n_64, n_60, in_0[1], in_0[0]);
  nand g5 (n_65, in_0[2], n_61, n_62);
  nand g6 (n_66, in_0[2], n_61, in_0[0]);
  nand g7 (n_67, in_0[2], in_0[1], n_62);
  nand g8 (n_39, in_0[2], in_0[1], in_0[0]);
  not g9 (out_0[7], n_25);
  not g10 (out_0[6], n_27);
  not g11 (out_0[5], n_63);
  not g12 (out_0[4], n_64);
  not g13 (out_0[3], n_65);
  not g14 (out_0[2], n_66);
  not g15 (out_0[1], n_67);
  not g16 (out_0[0], n_39);
  not g17 (n_60, in_0[2]);
  not g18 (n_61, in_0[1]);
  not g19 (n_62, in_0[0]);
endmodule

module fx68k_mux_1775(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [7:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [7:0] z;
  wire [7:0] ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [7:0] z;
  CDN_mux8 g1(.sel0 (ctl[7]), .data0 (in_0[7]), .sel1 (ctl[6]), .data1
       (in_1[7]), .sel2 (ctl[5]), .data2 (in_2[7]), .sel3 (ctl[4]),
       .data3 (in_3[7]), .sel4 (ctl[3]), .data4 (in_4[7]), .sel5
       (ctl[2]), .data5 (in_5[7]), .sel6 (ctl[1]), .data6 (in_6[7]),
       .sel7 (ctl[0]), .data7 (in_7[7]), .z (z[7]));
  CDN_mux8 g9(.sel0 (ctl[7]), .data0 (in_0[6]), .sel1 (ctl[6]), .data1
       (in_1[6]), .sel2 (ctl[5]), .data2 (in_2[6]), .sel3 (ctl[4]),
       .data3 (in_3[6]), .sel4 (ctl[3]), .data4 (in_4[6]), .sel5
       (ctl[2]), .data5 (in_5[6]), .sel6 (ctl[1]), .data6 (in_6[6]),
       .sel7 (ctl[0]), .data7 (in_7[6]), .z (z[6]));
  CDN_mux8 g10(.sel0 (ctl[7]), .data0 (in_0[5]), .sel1 (ctl[6]), .data1
       (in_1[5]), .sel2 (ctl[5]), .data2 (in_2[5]), .sel3 (ctl[4]),
       .data3 (in_3[5]), .sel4 (ctl[3]), .data4 (in_4[5]), .sel5
       (ctl[2]), .data5 (in_5[5]), .sel6 (ctl[1]), .data6 (in_6[5]),
       .sel7 (ctl[0]), .data7 (in_7[5]), .z (z[5]));
  CDN_mux8 g11(.sel0 (ctl[7]), .data0 (in_0[4]), .sel1 (ctl[6]), .data1
       (in_1[4]), .sel2 (ctl[5]), .data2 (in_2[4]), .sel3 (ctl[4]),
       .data3 (in_3[4]), .sel4 (ctl[3]), .data4 (in_4[4]), .sel5
       (ctl[2]), .data5 (in_5[4]), .sel6 (ctl[1]), .data6 (in_6[4]),
       .sel7 (ctl[0]), .data7 (in_7[4]), .z (z[4]));
  CDN_mux8 g12(.sel0 (ctl[7]), .data0 (in_0[3]), .sel1 (ctl[6]), .data1
       (in_1[3]), .sel2 (ctl[5]), .data2 (in_2[3]), .sel3 (ctl[4]),
       .data3 (in_3[3]), .sel4 (ctl[3]), .data4 (in_4[3]), .sel5
       (ctl[2]), .data5 (in_5[3]), .sel6 (ctl[1]), .data6 (in_6[3]),
       .sel7 (ctl[0]), .data7 (in_7[3]), .z (z[3]));
  CDN_mux8 g13(.sel0 (ctl[7]), .data0 (in_0[2]), .sel1 (ctl[6]), .data1
       (in_1[2]), .sel2 (ctl[5]), .data2 (in_2[2]), .sel3 (ctl[4]),
       .data3 (in_3[2]), .sel4 (ctl[3]), .data4 (in_4[2]), .sel5
       (ctl[2]), .data5 (in_5[2]), .sel6 (ctl[1]), .data6 (in_6[2]),
       .sel7 (ctl[0]), .data7 (in_7[2]), .z (z[2]));
  CDN_mux8 g14(.sel0 (ctl[7]), .data0 (in_0[1]), .sel1 (ctl[6]), .data1
       (in_1[1]), .sel2 (ctl[5]), .data2 (in_2[1]), .sel3 (ctl[4]),
       .data3 (in_3[1]), .sel4 (ctl[3]), .data4 (in_4[1]), .sel5
       (ctl[2]), .data5 (in_5[1]), .sel6 (ctl[1]), .data6 (in_6[1]),
       .sel7 (ctl[0]), .data7 (in_7[1]), .z (z[1]));
  CDN_mux8 g15(.sel0 (ctl[7]), .data0 (in_0[0]), .sel1 (ctl[6]), .data1
       (in_1[0]), .sel2 (ctl[5]), .data2 (in_2[0]), .sel3 (ctl[4]),
       .data3 (in_3[0]), .sel4 (ctl[3]), .data4 (in_4[0]), .sel5
       (ctl[2]), .data5 (in_5[0]), .sel6 (ctl[1]), .data6 (in_6[0]),
       .sel7 (ctl[0]), .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_bmux_1782(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, z);
  input [3:0] ctl;
  input [14:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15;
  output [14:0] z;
  wire [3:0] ctl;
  wire [14:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15;
  wire [14:0] z;
  CDN_bmux16 g1(.sel0 (ctl[0]), .data0 (in_0[14]), .data1 (in_1[14]),
       .sel1 (ctl[1]), .data2 (in_2[14]), .data3 (in_3[14]), .sel2
       (ctl[2]), .data4 (in_4[14]), .data5 (in_5[14]), .data6
       (in_6[14]), .data7 (in_7[14]), .sel3 (ctl[3]), .data8
       (in_8[14]), .data9 (in_9[14]), .data10 (in_10[14]), .data11
       (in_11[14]), .data12 (in_12[14]), .data13 (in_13[14]), .data14
       (in_14[14]), .data15 (in_15[14]), .z (z[14]));
  CDN_bmux16 g2(.sel0 (ctl[0]), .data0 (in_0[13]), .data1 (in_1[13]),
       .sel1 (ctl[1]), .data2 (in_2[13]), .data3 (in_3[13]), .sel2
       (ctl[2]), .data4 (in_4[13]), .data5 (in_5[13]), .data6
       (in_6[13]), .data7 (in_7[13]), .sel3 (ctl[3]), .data8
       (in_8[13]), .data9 (in_9[13]), .data10 (in_10[13]), .data11
       (in_11[13]), .data12 (in_12[13]), .data13 (in_13[13]), .data14
       (in_14[13]), .data15 (in_15[13]), .z (z[13]));
  CDN_bmux16 g3(.sel0 (ctl[0]), .data0 (in_0[12]), .data1 (in_1[12]),
       .sel1 (ctl[1]), .data2 (in_2[12]), .data3 (in_3[12]), .sel2
       (ctl[2]), .data4 (in_4[12]), .data5 (in_5[12]), .data6
       (in_6[12]), .data7 (in_7[12]), .sel3 (ctl[3]), .data8
       (in_8[12]), .data9 (in_9[12]), .data10 (in_10[12]), .data11
       (in_11[12]), .data12 (in_12[12]), .data13 (in_13[12]), .data14
       (in_14[12]), .data15 (in_15[12]), .z (z[12]));
  CDN_bmux16 g4(.sel0 (ctl[0]), .data0 (in_0[11]), .data1 (in_1[11]),
       .sel1 (ctl[1]), .data2 (in_2[11]), .data3 (in_3[11]), .sel2
       (ctl[2]), .data4 (in_4[11]), .data5 (in_5[11]), .data6
       (in_6[11]), .data7 (in_7[11]), .sel3 (ctl[3]), .data8
       (in_8[11]), .data9 (in_9[11]), .data10 (in_10[11]), .data11
       (in_11[11]), .data12 (in_12[11]), .data13 (in_13[11]), .data14
       (in_14[11]), .data15 (in_15[11]), .z (z[11]));
  CDN_bmux16 g5(.sel0 (ctl[0]), .data0 (in_0[10]), .data1 (in_1[10]),
       .sel1 (ctl[1]), .data2 (in_2[10]), .data3 (in_3[10]), .sel2
       (ctl[2]), .data4 (in_4[10]), .data5 (in_5[10]), .data6
       (in_6[10]), .data7 (in_7[10]), .sel3 (ctl[3]), .data8
       (in_8[10]), .data9 (in_9[10]), .data10 (in_10[10]), .data11
       (in_11[10]), .data12 (in_12[10]), .data13 (in_13[10]), .data14
       (in_14[10]), .data15 (in_15[10]), .z (z[10]));
  CDN_bmux16 g6(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .sel2
       (ctl[2]), .data4 (in_4[9]), .data5 (in_5[9]), .data6 (in_6[9]),
       .data7 (in_7[9]), .sel3 (ctl[3]), .data8 (in_8[9]), .data9
       (in_9[9]), .data10 (in_10[9]), .data11 (in_11[9]), .data12
       (in_12[9]), .data13 (in_13[9]), .data14 (in_14[9]), .data15
       (in_15[9]), .z (z[9]));
  CDN_bmux16 g7(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .sel2
       (ctl[2]), .data4 (in_4[8]), .data5 (in_5[8]), .data6 (in_6[8]),
       .data7 (in_7[8]), .sel3 (ctl[3]), .data8 (in_8[8]), .data9
       (in_9[8]), .data10 (in_10[8]), .data11 (in_11[8]), .data12
       (in_12[8]), .data13 (in_13[8]), .data14 (in_14[8]), .data15
       (in_15[8]), .z (z[8]));
  CDN_bmux16 g8(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .data7 (in_7[7]), .sel3 (ctl[3]), .data8 (in_8[7]), .data9
       (in_9[7]), .data10 (in_10[7]), .data11 (in_11[7]), .data12
       (in_12[7]), .data13 (in_13[7]), .data14 (in_14[7]), .data15
       (in_15[7]), .z (z[7]));
  CDN_bmux16 g9(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .data7 (in_7[6]), .sel3 (ctl[3]), .data8 (in_8[6]), .data9
       (in_9[6]), .data10 (in_10[6]), .data11 (in_11[6]), .data12
       (in_12[6]), .data13 (in_13[6]), .data14 (in_14[6]), .data15
       (in_15[6]), .z (z[6]));
  CDN_bmux16 g10(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .data7 (in_7[5]), .sel3 (ctl[3]), .data8 (in_8[5]), .data9
       (in_9[5]), .data10 (in_10[5]), .data11 (in_11[5]), .data12
       (in_12[5]), .data13 (in_13[5]), .data14 (in_14[5]), .data15
       (in_15[5]), .z (z[5]));
  CDN_bmux16 g11(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .data7 (in_7[4]), .sel3 (ctl[3]), .data8 (in_8[4]), .data9
       (in_9[4]), .data10 (in_10[4]), .data11 (in_11[4]), .data12
       (in_12[4]), .data13 (in_13[4]), .data14 (in_14[4]), .data15
       (in_15[4]), .z (z[4]));
  CDN_bmux16 g12(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .sel3 (ctl[3]), .data8 (in_8[3]), .data9
       (in_9[3]), .data10 (in_10[3]), .data11 (in_11[3]), .data12
       (in_12[3]), .data13 (in_13[3]), .data14 (in_14[3]), .data15
       (in_15[3]), .z (z[3]));
  CDN_bmux16 g13(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .sel3 (ctl[3]), .data8 (in_8[2]), .data9
       (in_9[2]), .data10 (in_10[2]), .data11 (in_11[2]), .data12
       (in_12[2]), .data13 (in_13[2]), .data14 (in_14[2]), .data15
       (in_15[2]), .z (z[2]));
  CDN_bmux16 g14(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .sel3 (ctl[3]), .data8 (in_8[1]), .data9
       (in_9[1]), .data10 (in_10[1]), .data11 (in_11[1]), .data12
       (in_12[1]), .data13 (in_13[1]), .data14 (in_14[1]), .data15
       (in_15[1]), .z (z[1]));
  CDN_bmux16 g15(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .sel3 (ctl[3]), .data8 (in_8[0]), .data9
       (in_9[0]), .data10 (in_10[0]), .data11 (in_11[0]), .data12
       (in_12[0]), .data13 (in_13[0]), .data14 (in_14[0]), .data15
       (in_15[0]), .z (z[0]));
endmodule

module fx68k_mux_1783(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input in_0, in_1;
  output z;
  wire [1:0] ctl;
  wire in_0, in_1;
  wire z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0), .sel1 (ctl[0]), .data1
       (in_1), .z (z));
endmodule

module fx68k_rowDecoder(ird, row, noCcrEn, isArX);
  input [15:0] ird;
  output [15:0] row;
  output noCcrEn, isArX;
  wire [15:0] ird;
  wire [15:0] row;
  wire noCcrEn, isArX;
  wire [1:0] stype;
  wire _X_, eaAdir, eaRdir, n_6, n_7, n_8, n_9, n_11;
  wire n_13, n_22, n_32, n_782, n_783, n_784, n_785, n_786;
  wire n_787, n_788, n_790, n_792, n_793, n_794, n_795, n_796;
  wire n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804;
  wire n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_817, n_818, n_819, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837;
  wire n_838, n_839, n_841, n_842, n_844, n_846, n_847, n_853;
  wire n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_865;
  wire n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_908;
  wire n_909, n_912, n_918, n_919, n_920, n_926, n_927, n_944;
  wire n_945, n_946, n_947, n_954, n_958, n_959, n_960, n_963;
  wire size11;
  assign row[0] = 1'b0;
  fx68k_case_box_1045 ctl_ird_650_16(.in_0 (ird[11:9]), .out_0 ({n_782,
       n_783, n_784, n_785, n_786, n_787, n_788}));
  fx68k_mux_1738 mux_row_650_16(.ctl ({n_782, n_783, n_784, n_785,
       n_786, n_787, n_788}), .in_0 (6'b000100), .in_1 (6'b000001),
       .in_2 (6'b000010), .in_3 (6'b001000), .in_4 ({1'b1, _X_, _X_,
       _X_, _X_, _X_}), .in_5 (6'b010000), .in_6 (6'b000000), .z
       ({n_790, n_799, n_798, n_797, n_794, n_793}));
  fx68k_bmux_1520 mux_655_20(.ctl (ird[7]), .in_0 (2'b10), .in_1
       (2'b01), .z ({n_796, n_795}));
  fx68k_mux_1744 mux_row_650_29(.ctl ({n_790, n_792}), .in_0 ({3'b000,
       n_796, n_795, 2'b00}), .in_1 ({n_799, n_798, n_797, 2'b00,
       n_794, n_793}), .z ({n_806, n_805, n_804, n_803, n_802, n_801,
       n_800}));
  fx68k_bmux mux_row_648_9(.ctl (ird[8]), .in_0 ({n_806, n_805, n_804,
       n_803, n_802, 1'b0, n_801, n_800}), .in_1 (8'b00000100), .z
       ({n_900, n_893, n_890, n_887, n_885, n_881, n_876, n_872}));
  fx68k_bmux_1520 mux_663_12(.ctl (ird[7]), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_832, n_830}));
  fx68k_case_box_1049 ctl_ird_664_16(.in_0 (ird[11:9]), .out_0 ({n_807,
       n_808, n_809, n_810, n_811, n_812, n_813, n_814}));
  fx68k_mux_893 mux_row_664_16(.ctl ({n_807, n_808, n_809, n_810,
       n_811, n_812, n_813, n_814}), .in_0 (7'b0100000), .in_1
       (7'b0000010), .in_2 (7'b0000100), .in_3 (7'b0000001), .in_4
       ({1'b1, _X_, _X_, _X_, _X_, _X_, _X_}), .in_5 (7'b0010000),
       .in_6 (7'b0001000), .in_7 (7'b0000000), .z ({n_815, n_825,
       n_823, n_821, n_820, n_819, n_818}));
  fx68k_bmux_1520 mux_669_21(.ctl (ird[7]), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_824, n_822}));
  fx68k_mux_1759 mux_row_664_30(.ctl ({n_815, n_817}), .in_0 ({n_824,
       n_822, 4'b0000}), .in_1 ({n_825, n_823, n_821, n_820, n_819,
       n_818}), .z ({n_833, n_831, n_829, n_828, n_827, n_826}));
  fx68k_bmux_1505 mux_row_662_9(.ctl (ird[8]), .in_0 ({n_833, n_831,
       n_829, n_828, n_827, n_826}), .in_1 ({n_832, n_830, 4'b0000}),
       .z ({n_898, n_896, n_882, n_877, n_873, n_866}));
  fx68k_bmux_1520 mux_686_11(.ctl (ird[8]), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_835, n_834}));
  fx68k_bmux_1766 mux_row_683_8(.ctl (size11), .in_0 ({1'b0, n_835,
       n_834}), .in_1 (3'b100), .z ({n_901, n_878, n_867}));
  fx68k_bmux_1520 mux_row_692_20(.ctl (n_836), .in_0 (2'b10), .in_1
       (2'b01), .z ({n_838, n_837}));
  fx68k_bmux_1766 mux_row_690_8(.ctl (size11), .in_0 ({n_838, n_837,
       1'b0}), .in_1 (3'b001), .z ({n_899, n_888, n_865}));
  fx68k_mux_1769 mux_row_697_25(.ctl ({n_839, n_841}), .in_0 (2'b10),
       .in_1 (2'b01), .z ({n_891, n_879}));
  fx68k_mux_1769 mux_row_702_25(.ctl ({n_842, n_844}), .in_0 (2'b10),
       .in_1 (2'b01), .z ({n_897, n_883}));
  fx68k_bmux_1520 mux_row_709_20(.ctl (n_836), .in_0 (2'b10), .in_1
       (2'b01), .z ({n_847, n_846}));
  fx68k_bmux_1766 mux_row_707_8(.ctl (size11), .in_0 ({1'b0, n_847,
       n_846}), .in_1 (3'b100), .z ({n_884, n_874, n_870}));
  fx68k_mux_1769 mux_row_714_25(.ctl ({n_839, n_841}), .in_0 (2'b10),
       .in_1 (2'b01), .z ({n_895, n_868}));
  fx68k_bmux_1520 mux_stype_722_9(.ctl (size11), .in_0 (ird[4:3]),
       .in_1 (ird[10:9]), .z (stype));
  fx68k_case_box_1064 ctl_727_5(.in_0 ({stype, ird[8]}), .out_0
       ({n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860}));
  fx68k_mux_1775 mux_row_727_5(.ctl ({n_853, n_854, n_855, n_856,
       n_857, n_858, n_859, n_860}), .in_0 (8'b00000001), .in_1
       (8'b00000010), .in_2 (8'b00001000), .in_3 (8'b00000100), .in_4
       (8'b00010000), .in_5 (8'b10000000), .in_6 (8'b01000000), .in_7
       (8'b00100000), .z ({n_894, n_892, n_889, n_886, n_880, n_875,
       n_871, n_869}));
  fx68k_bmux_1782 mux_row_645_16(.ctl (ird[15:12]), .in_0 ({1'b0,
       n_898, n_896, 6'b000000, n_882, n_877, n_873, 1'b0, n_866,
       1'b0}), .in_1 (15'b000000000000010), .in_2
       (15'b000000000000010), .in_3 (15'b000000000000010), .in_4
       ({n_900, 3'b000, n_893, n_890, n_887, n_885, 1'b0, n_881, n_876,
       n_872, 3'b000}), .in_5 ({n_901, 9'b000000000, n_878, 2'b00,
       n_867, 1'b0}), .in_6 (15'b000000000000000), .in_7
       (15'b000000000000010), .in_8 ({1'b0, n_899, 4'b0000, n_888,
       7'b0000000, n_865}), .in_9 ({5'b00000, n_891, 4'b0000, n_879,
       4'b0000}), .in_10 (15'b000000000000000), .in_11 ({2'b00, n_897,
       6'b000000, n_883, 5'b00000}), .in_12 ({8'b00000000, n_884,
       2'b00, n_874, n_870, 2'b00}), .in_13 ({3'b000, n_895,
       9'b000000000, n_868, 1'b0}), .in_14 ({4'b0000, n_894, n_892,
       n_889, n_886, 2'b00, n_880, n_875, n_871, n_869, 1'b0}), .in_15
       (15'b000000000000000), .z (row[15:1]));
  fx68k_mux_1783 mux_isArX_634_9(.ctl ({n_902, n_903}), .in_0 (n_904),
       .in_1 (1'b0), .z (isArX));
  and g1 (size11, ird[7], ird[6]);
  or g2 (n_904, row[10], row[12]);
  and g3 (n_836, ird[8], eaRdir);
  not g4 (n_908, size11);
  and g5 (n_909, ird[8], n_908);
  and g6 (n_839, n_909, eaRdir);
  and g10 (n_842, n_909, n_912);
  not g15 (n_22, ird[13]);
  and g19 (n_920, n_918, eaAdir);
  or g20 (n_926, n_919, n_920);
  or g26 (noCcrEn, n_926, n_927);
  CDN_dc logicX_inst(.cf (1'b0), .dcf (1'b1), .z (_X_));
  not g35 (n_945, ird[5]);
  nand g36 (n_946, n_944, n_945);
  not g37 (eaRdir, n_946);
  nor g39 (n_947, ird[5], ird[4]);
  nand g40 (n_912, n_947, ird[3]);
  not g41 (eaAdir, n_912);
  not g45 (n_6, ird[15]);
  nand g46 (n_954, n_6, ird[12], n_22, ird[14]);
  not g47 (n_918, n_954);
  not g52 (n_944, ird[4]);
  and g53 (n_919, ird[15], n_22, ird[12], size11);
  nor g54 (n_959, ird[14], ird[8]);
  and g55 (n_960, n_958, n_6);
  not g56 (n_958, ird[7]);
  and g57 (n_927, ird[13], ird[6], n_959, n_960);
  not g58 (n_792, n_790);
  not g61 (n_817, n_815);
  not g65 (n_841, n_839);
  not g67 (n_844, n_842);
  not g70 (n_903, n_902);
  nor g18 (n_902, ird[13], n_13);
  nand g73 (n_13, n_9, n_32);
  not g74 (n_963, ird[12]);
  and g75 (n_7, ird[12], ird[15]);
  and g7 (n_8, n_963, n_6);
  or g8 (n_9, n_7, n_8);
  nand g9 (n_32, n_6, n_11);
  not g77 (n_11, ird[14]);
endmodule

module fx68k_case_box_1075(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_mux_1788(ctl, in_0, in_1, in_2, z);
  input [2:0] ctl;
  input [4:0] in_0, in_1, in_2;
  output [4:0] z;
  wire [2:0] ctl;
  wire [4:0] in_0, in_1, in_2;
  wire [4:0] z;
  CDN_mux3 g1(.sel0 (ctl[2]), .data0 (in_0[4]), .sel1 (ctl[1]), .data1
       (in_1[4]), .sel2 (ctl[0]), .data2 (in_2[4]), .z (z[4]));
  CDN_mux3 g6(.sel0 (ctl[2]), .data0 (in_0[3]), .sel1 (ctl[1]), .data1
       (in_1[3]), .sel2 (ctl[0]), .data2 (in_2[3]), .z (z[3]));
  CDN_mux3 g7(.sel0 (ctl[2]), .data0 (in_0[2]), .sel1 (ctl[1]), .data1
       (in_1[2]), .sel2 (ctl[0]), .data2 (in_2[2]), .z (z[2]));
  CDN_mux3 g8(.sel0 (ctl[2]), .data0 (in_0[1]), .sel1 (ctl[1]), .data1
       (in_1[1]), .sel2 (ctl[0]), .data2 (in_2[1]), .z (z[1]));
  CDN_mux3 g9(.sel0 (ctl[2]), .data0 (in_0[0]), .sel1 (ctl[1]), .data1
       (in_1[0]), .sel2 (ctl[0]), .data2 (in_2[0]), .z (z[0]));
endmodule

module fx68k_case_box_1076(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_mux_1792(ctl, in_0, in_1, in_2, z);
  input [2:0] ctl;
  input [3:0] in_0, in_1, in_2;
  output [3:0] z;
  wire [2:0] ctl;
  wire [3:0] in_0, in_1, in_2;
  wire [3:0] z;
  CDN_mux3 g1(.sel0 (ctl[2]), .data0 (in_0[3]), .sel1 (ctl[1]), .data1
       (in_1[3]), .sel2 (ctl[0]), .data2 (in_2[3]), .z (z[3]));
  CDN_mux3 g5(.sel0 (ctl[2]), .data0 (in_0[2]), .sel1 (ctl[1]), .data1
       (in_1[2]), .sel2 (ctl[0]), .data2 (in_2[2]), .z (z[2]));
  CDN_mux3 g6(.sel0 (ctl[2]), .data0 (in_0[1]), .sel1 (ctl[1]), .data1
       (in_1[1]), .sel2 (ctl[0]), .data2 (in_2[1]), .z (z[1]));
  CDN_mux3 g7(.sel0 (ctl[2]), .data0 (in_0[0]), .sel1 (ctl[1]), .data1
       (in_1[0]), .sel2 (ctl[0]), .data2 (in_2[0]), .z (z[0]));
endmodule

module fx68k_case_box_1082(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_mux_1800(ctl, in_0, in_1, in_2, z);
  input [2:0] ctl, in_0, in_1, in_2;
  output [2:0] z;
  wire [2:0] ctl, in_0, in_1, in_2;
  wire [2:0] z;
  CDN_mux3 g1(.sel0 (ctl[2]), .data0 (in_0[2]), .sel1 (ctl[1]), .data1
       (in_1[2]), .sel2 (ctl[0]), .data2 (in_2[2]), .z (z[2]));
  CDN_mux3 g4(.sel0 (ctl[2]), .data0 (in_0[1]), .sel1 (ctl[1]), .data1
       (in_1[1]), .sel2 (ctl[0]), .data2 (in_2[1]), .z (z[1]));
  CDN_mux3 g5(.sel0 (ctl[2]), .data0 (in_0[0]), .sel1 (ctl[1]), .data1
       (in_1[0]), .sel2 (ctl[0]), .data2 (in_2[0]), .z (z[0]));
endmodule

module fx68k_case_box_1085(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_case_box_1088(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_case_box_1091(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_case_box_1094(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_case_box_1097(in_0, out_0);
  input [2:0] in_0;
  output [3:0] out_0;
  wire [2:0] in_0;
  wire [3:0] out_0;
  assign out_0[0] = 1'b0;
  assign out_0[1] = in_0[2];
  assign out_0[2] = in_0[0];
  nor g1 (out_0[3], in_0[2], in_0[0]);
endmodule

module fx68k_mux_1814(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, in_13, z);
  input [13:0] ctl;
  input [4:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13;
  output [4:0] z;
  wire [13:0] ctl;
  wire [4:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13;
  wire [4:0] z;
  CDN_mux14 g1(.sel0 (ctl[13]), .data0 (in_0[4]), .sel1 (ctl[12]),
       .data1 (in_1[4]), .sel2 (ctl[11]), .data2 (in_2[4]), .sel3
       (ctl[10]), .data3 (in_3[4]), .sel4 (ctl[9]), .data4 (in_4[4]),
       .sel5 (ctl[8]), .data5 (in_5[4]), .sel6 (ctl[7]), .data6
       (in_6[4]), .sel7 (ctl[6]), .data7 (in_7[4]), .sel8 (ctl[5]),
       .data8 (in_8[4]), .sel9 (ctl[4]), .data9 (in_9[4]), .sel10
       (ctl[3]), .data10 (in_10[4]), .sel11 (ctl[2]), .data11
       (in_11[4]), .sel12 (ctl[1]), .data12 (in_12[4]), .sel13
       (ctl[0]), .data13 (in_13[4]), .z (z[4]));
  CDN_mux14 g6(.sel0 (ctl[13]), .data0 (in_0[3]), .sel1 (ctl[12]),
       .data1 (in_1[3]), .sel2 (ctl[11]), .data2 (in_2[3]), .sel3
       (ctl[10]), .data3 (in_3[3]), .sel4 (ctl[9]), .data4 (in_4[3]),
       .sel5 (ctl[8]), .data5 (in_5[3]), .sel6 (ctl[7]), .data6
       (in_6[3]), .sel7 (ctl[6]), .data7 (in_7[3]), .sel8 (ctl[5]),
       .data8 (in_8[3]), .sel9 (ctl[4]), .data9 (in_9[3]), .sel10
       (ctl[3]), .data10 (in_10[3]), .sel11 (ctl[2]), .data11
       (in_11[3]), .sel12 (ctl[1]), .data12 (in_12[3]), .sel13
       (ctl[0]), .data13 (in_13[3]), .z (z[3]));
  CDN_mux14 g7(.sel0 (ctl[13]), .data0 (in_0[2]), .sel1 (ctl[12]),
       .data1 (in_1[2]), .sel2 (ctl[11]), .data2 (in_2[2]), .sel3
       (ctl[10]), .data3 (in_3[2]), .sel4 (ctl[9]), .data4 (in_4[2]),
       .sel5 (ctl[8]), .data5 (in_5[2]), .sel6 (ctl[7]), .data6
       (in_6[2]), .sel7 (ctl[6]), .data7 (in_7[2]), .sel8 (ctl[5]),
       .data8 (in_8[2]), .sel9 (ctl[4]), .data9 (in_9[2]), .sel10
       (ctl[3]), .data10 (in_10[2]), .sel11 (ctl[2]), .data11
       (in_11[2]), .sel12 (ctl[1]), .data12 (in_12[2]), .sel13
       (ctl[0]), .data13 (in_13[2]), .z (z[2]));
  CDN_mux14 g8(.sel0 (ctl[13]), .data0 (in_0[1]), .sel1 (ctl[12]),
       .data1 (in_1[1]), .sel2 (ctl[11]), .data2 (in_2[1]), .sel3
       (ctl[10]), .data3 (in_3[1]), .sel4 (ctl[9]), .data4 (in_4[1]),
       .sel5 (ctl[8]), .data5 (in_5[1]), .sel6 (ctl[7]), .data6
       (in_6[1]), .sel7 (ctl[6]), .data7 (in_7[1]), .sel8 (ctl[5]),
       .data8 (in_8[1]), .sel9 (ctl[4]), .data9 (in_9[1]), .sel10
       (ctl[3]), .data10 (in_10[1]), .sel11 (ctl[2]), .data11
       (in_11[1]), .sel12 (ctl[1]), .data12 (in_12[1]), .sel13
       (ctl[0]), .data13 (in_13[1]), .z (z[1]));
  CDN_mux14 g9(.sel0 (ctl[13]), .data0 (in_0[0]), .sel1 (ctl[12]),
       .data1 (in_1[0]), .sel2 (ctl[11]), .data2 (in_2[0]), .sel3
       (ctl[10]), .data3 (in_3[0]), .sel4 (ctl[9]), .data4 (in_4[0]),
       .sel5 (ctl[8]), .data5 (in_5[0]), .sel6 (ctl[7]), .data6
       (in_6[0]), .sel7 (ctl[6]), .data7 (in_7[0]), .sel8 (ctl[5]),
       .data8 (in_8[0]), .sel9 (ctl[4]), .data9 (in_9[0]), .sel10
       (ctl[3]), .data10 (in_10[0]), .sel11 (ctl[2]), .data11
       (in_11[0]), .sel12 (ctl[1]), .data12 (in_12[0]), .sel13
       (ctl[0]), .data13 (in_13[0]), .z (z[0]));
endmodule

module fx68k_aluGetOp(row, col, isCorf, aluOp);
  input [15:0] row;
  input [2:0] col;
  input isCorf;
  output [4:0] aluOp;
  wire [15:0] row;
  wire [2:0] col;
  wire isCorf;
  wire [4:0] aluOp;
  wire UNCONNECTED428, UNCONNECTED429, UNCONNECTED430, UNCONNECTED431,
       UNCONNECTED432, UNCONNECTED433, UNCONNECTED434, UNCONNECTED435;
  wire n_6, n_8, n_62, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_207, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_251, n_261, n_262, n_263, n_264, n_265, n_266, n_267;
  wire n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275;
  wire n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283;
  wire n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291;
  wire n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299;
  wire n_300, n_301, n_302, n_303, n_304, n_305, n_311, n_314;
  wire n_318;
  fx68k_case_box_1075 ctl_col_538_19(.in_0 (col), .out_0 ({n_200,
       n_201, n_202, UNCONNECTED428}));
  fx68k_mux_1788 mux_aluOp_538_19(.ctl ({n_200, n_201, n_202}), .in_0
       (5'b00010), .in_1 (5'b01010), .in_2 (5'b10101), .z ({n_290,
       n_283, n_275, n_268, n_261}));
  fx68k_case_box_1076 ctl_col_545_19(.in_0 (col), .out_0 ({n_203,
       n_204, n_205, UNCONNECTED429}));
  fx68k_mux_1792 mux_aluOp_545_19(.ctl ({n_203, n_204, n_205}), .in_0
       (4'b0100), .in_1 (4'b1011), .in_2 (4'b1110), .z ({n_284, n_276,
       n_269, n_262}));
  fx68k_bmux_1520 mux_554_17(.ctl (isCorf), .in_0 (2'b00), .in_1
       (2'b11), .z ({n_211, n_210}));
  fx68k_mux_1792 mux_aluOp_552_19(.ctl ({n_207, col[0], col[2]}), .in_0
       (4'b0100), .in_1 ({n_211, 1'b0, n_210, 1'b0}), .in_2 (4'b0101),
       .z ({n_291, n_285, n_270, n_263}));
  fx68k_bmux_1766 mux_559_20(.ctl (n_212), .in_0 (3'b000), .in_1
       (3'b111), .z ({n_286, n_277, n_271}));
  fx68k_case_box_1082 ctl_col_563_19(.in_0 (col), .out_0 ({n_213,
       n_214, n_215, UNCONNECTED430}));
  fx68k_mux_1800 mux_aluOp_563_19(.ctl ({n_213, n_214, n_215}), .in_0
       (3'b001), .in_1 (3'b011), .in_2 (3'b100), .z ({n_292, n_287,
       n_272}));
  fx68k_case_box_1085 ctl_col_570_19(.in_0 (col), .out_0 ({n_216,
       n_217, n_218, UNCONNECTED431}));
  fx68k_mux_1800 mux_aluOp_570_19(.ctl ({n_216, n_217, n_218}), .in_0
       (3'b001), .in_1 (3'b010), .in_2 (3'b110), .z ({n_293, n_278,
       n_273}));
  fx68k_case_box_1088 ctl_col_579_19(.in_0 (col), .out_0 ({n_219,
       n_220, n_221, UNCONNECTED432}));
  fx68k_mux_1800 mux_aluOp_579_19(.ctl ({n_219, n_220, n_221}), .in_0
       (3'b011), .in_1 (3'b001), .in_2 (3'b110), .z ({n_294, n_279,
       n_264}));
  fx68k_case_box_1091 ctl_col_586_19(.in_0 (col), .out_0 ({n_222,
       n_223, n_224, UNCONNECTED433}));
  fx68k_mux_1792 mux_aluOp_586_19(.ctl ({n_222, n_223, n_224}), .in_0
       (4'b0011), .in_1 (4'b0110), .in_2 (4'b1001), .z ({n_295, n_280,
       n_274, n_265}));
  fx68k_case_box_1094 ctl_col_593_19(.in_0 (col), .out_0 ({n_225,
       n_226, n_227, UNCONNECTED434}));
  fx68k_mux_1800 mux_aluOp_593_19(.ctl ({n_225, n_226, n_227}), .in_0
       (3'b001), .in_1 (3'b010), .in_2 (3'b100), .z ({n_296, n_288,
       n_266}));
  fx68k_case_box_1097 ctl_col_600_19(.in_0 (col), .out_0 ({n_228,
       n_229, n_230, UNCONNECTED435}));
  fx68k_mux_1694 mux_aluOp_600_19(.ctl ({n_228, n_229, n_230}), .in_0
       (2'b01), .in_1 (2'b01), .in_2 (2'b10), .z ({n_297, n_281}));
  fx68k_bmux_1503 mux_608_27(.ctl (n_212), .in_0 (1'b0), .in_1 (1'b1),
       .z (n_267));
  fx68k_bmux_1520 mux_609_27(.ctl (n_231), .in_0 (2'b10), .in_1
       (2'b01), .z ({n_289, n_282}));
  fx68k_mux_1814 mux_aluOp_536_11(.ctl ({row[1], row[2], row[3],
       row[4], n_251, row[7], row[8], row[9], row[10], row[11],
       row[12], row[13], row[14], row[15]}), .in_0 ({n_290, n_283,
       n_275, n_268, n_261}), .in_1 ({1'b0, n_284, n_276, n_269,
       n_262}), .in_2 ({n_291, n_285, 1'b1, n_270, n_263}), .in_3
       ({1'b0, n_286, n_277, n_271, 1'b1}), .in_4 ({n_292, n_287, 1'b0,
       n_272, 1'b0}), .in_5 ({n_293, 1'b0, n_278, n_273, 1'b0}), .in_6
       ({n_294, 1'b0, n_279, 1'b0, n_264}), .in_7 ({n_295, 1'b0, n_280,
       n_274, n_265}), .in_8 ({n_296, n_288, 2'b01, n_266}), .in_9
       ({n_297, 1'b0, n_281, 2'b11}), .in_10 (5'b01100), .in_11
       (5'b01001), .in_12 ({4'b0100, n_267}), .in_13 ({1'b0, n_289,
       n_282, 2'b00}), .z ({n_305, n_304, n_303, n_302, n_301}));
  fx68k_mux_1788 mux_aluOp_531_16(.ctl ({n_298, n_299, n_300}), .in_0
       (5'b00001), .in_1 (5'b00101), .in_2 ({n_305, n_304, n_303,
       n_302, n_301}), .z (aluOp));
  nand g7 (n_314, n_311, n_8, col[2]);
  not g8 (n_212, n_314);
  not g11 (n_6, col[2]);
  nand g12 (n_318, n_6, col[0], col[1]);
  not g13 (n_231, n_318);
  not g14 (n_311, col[0]);
  not g15 (n_8, col[1]);
  nor g1 (n_207, col[2], col[0]);
  nor g27 (n_62, row[6], row[5]);
  not g28 (n_251, n_62);
  nor g37 (n_298, col[2], n_300);
  nand g38 (n_300, n_8, col[0]);
  nor g39 (n_299, n_300, n_6);
endmodule

module fx68k_mux_1828(ctl, in_0, in_1, in_2, in_3, in_4, in_5, z);
  input [5:0] ctl;
  input [4:0] in_0, in_1, in_2, in_3, in_4, in_5;
  output [4:0] z;
  wire [5:0] ctl;
  wire [4:0] in_0, in_1, in_2, in_3, in_4, in_5;
  wire [4:0] z;
  CDN_mux6 g1(.sel0 (ctl[5]), .data0 (in_0[4]), .sel1 (ctl[4]), .data1
       (in_1[4]), .sel2 (ctl[3]), .data2 (in_2[4]), .sel3 (ctl[2]),
       .data3 (in_3[4]), .sel4 (ctl[1]), .data4 (in_4[4]), .sel5
       (ctl[0]), .data5 (in_5[4]), .z (z[4]));
  CDN_mux6 g6(.sel0 (ctl[5]), .data0 (in_0[3]), .sel1 (ctl[4]), .data1
       (in_1[3]), .sel2 (ctl[3]), .data2 (in_2[3]), .sel3 (ctl[2]),
       .data3 (in_3[3]), .sel4 (ctl[1]), .data4 (in_4[3]), .sel5
       (ctl[0]), .data5 (in_5[3]), .z (z[3]));
  CDN_mux6 g7(.sel0 (ctl[5]), .data0 (in_0[2]), .sel1 (ctl[4]), .data1
       (in_1[2]), .sel2 (ctl[3]), .data2 (in_2[2]), .sel3 (ctl[2]),
       .data3 (in_3[2]), .sel4 (ctl[1]), .data4 (in_4[2]), .sel5
       (ctl[0]), .data5 (in_5[2]), .z (z[2]));
  CDN_mux6 g8(.sel0 (ctl[5]), .data0 (in_0[1]), .sel1 (ctl[4]), .data1
       (in_1[1]), .sel2 (ctl[3]), .data2 (in_2[1]), .sel3 (ctl[2]),
       .data3 (in_3[1]), .sel4 (ctl[1]), .data4 (in_4[1]), .sel5
       (ctl[0]), .data5 (in_5[1]), .z (z[1]));
  CDN_mux6 g9(.sel0 (ctl[5]), .data0 (in_0[0]), .sel1 (ctl[4]), .data1
       (in_1[0]), .sel2 (ctl[3]), .data2 (in_2[0]), .sel3 (ctl[2]),
       .data3 (in_3[0]), .sel4 (ctl[1]), .data4 (in_4[0]), .sel5
       (ctl[0]), .data5 (in_5[0]), .z (z[0]));
endmodule

module fx68k_case_box_1117(in_0, out_0);
  input [15:0] in_0;
  output [4:0] out_0;
  wire [15:0] in_0;
  wire [4:0] out_0;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  assign out_0[0] = 1'b0;
  assign out_0[3] = in_0[7];
  nor g1 (out_0[4], n_312, n_315);
  nand g2 (n_312, n_310, n_311);
  not g3 (n_310, in_0[7]);
  not g4 (n_311, in_0[10]);
  nand g5 (n_315, n_313, n_314);
  not g6 (n_313, in_0[11]);
  nor g7 (n_314, in_0[8], in_0[9]);
  nand g8 (out_0[2], n_311, n_316);
  not g9 (n_316, in_0[9]);
  nand g10 (out_0[1], n_313, n_317);
  not g11 (n_317, in_0[8]);
endmodule

module fx68k_mux_1834(ctl, in_0, in_1, in_2, in_3, z);
  input [3:0] ctl;
  input [4:0] in_0, in_1, in_2, in_3;
  output [4:0] z;
  wire [3:0] ctl;
  wire [4:0] in_0, in_1, in_2, in_3;
  wire [4:0] z;
  CDN_mux4 g1(.sel0 (ctl[3]), .data0 (in_0[4]), .sel1 (ctl[2]), .data1
       (in_1[4]), .sel2 (ctl[1]), .data2 (in_2[4]), .sel3 (ctl[0]),
       .data3 (in_3[4]), .z (z[4]));
  CDN_mux4 g6(.sel0 (ctl[3]), .data0 (in_0[3]), .sel1 (ctl[2]), .data1
       (in_1[3]), .sel2 (ctl[1]), .data2 (in_2[3]), .sel3 (ctl[0]),
       .data3 (in_3[3]), .z (z[3]));
  CDN_mux4 g7(.sel0 (ctl[3]), .data0 (in_0[2]), .sel1 (ctl[2]), .data1
       (in_1[2]), .sel2 (ctl[1]), .data2 (in_2[2]), .sel3 (ctl[0]),
       .data3 (in_3[2]), .z (z[2]));
  CDN_mux4 g8(.sel0 (ctl[3]), .data0 (in_0[1]), .sel1 (ctl[2]), .data1
       (in_1[1]), .sel2 (ctl[1]), .data2 (in_2[1]), .sel3 (ctl[0]),
       .data3 (in_3[1]), .z (z[1]));
  CDN_mux4 g9(.sel0 (ctl[3]), .data0 (in_0[0]), .sel1 (ctl[2]), .data1
       (in_1[0]), .sel2 (ctl[1]), .data2 (in_2[0]), .sel3 (ctl[0]),
       .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_ccrTable(col, row, finish, ccrMask);
  input [2:0] col;
  input [15:0] row;
  input finish;
  output [4:0] ccrMask;
  wire [2:0] col;
  wire [15:0] row;
  wire finish;
  wire [4:0] ccrMask;
  wire [4:0] ccrMask1;
  wire UNCONNECTED436, n_4, n_7, n_43, n_44, n_45, n_46, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_113, n_114;
  wire n_115, n_116, n_118, n_120, n_121, n_122, n_123, n_127;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_149;
  fx68k_bmux_1520 mux_833_15(.ctl (row[7]), .in_0 (2'b00), .in_1
       (2'b11), .z ({n_94, n_92}));
  fx68k_bmux_1766 mux_835_23(.ctl (n_91), .in_0 (3'b111), .in_1
       (3'b000), .z ({n_96, n_95, n_93}));
  fx68k_bmux_1766 mux_ccrMask1_832_7(.ctl (finish), .in_0 ({n_96, n_95,
       n_93}), .in_1 ({1'b1, n_94, n_92}), .z ({ccrMask1[3],
       ccrMask1[1:0]}));
  fx68k_bmux_1503 mux_789_22(.ctl (n_97), .in_0 (1'b1), .in_1 (1'b0),
       .z (n_118));
  fx68k_mux_1828 mux_ccrMask_784_11(.ctl ({row[1], n_113, n_114, n_115,
       n_116, row[15]}), .in_0 (5'b01111), .in_1 ({2'b11, n_118,
       2'b11}), .in_2 (5'b11111), .in_3 (5'b01111), .in_4 (5'b01111),
       .in_5 (5'b00000), .z ({n_139, n_137, n_135, n_133, n_131}));
  fx68k_case_box_1117 ctl_row_808_17(.in_0 (row), .out_0 ({n_120,
       n_121, n_122, n_123, UNCONNECTED436}));
  fx68k_mux_1577 mux_ccrMask_808_17(.ctl ({n_120, n_121, n_122,
       n_123}), .in_0 (1'b1), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b1),
       .z (n_140));
  fx68k_bmux_1504 mux_825_18(.ctl (row[1]), .in_0 (4'b0000), .in_1
       (4'b1111), .z ({n_138, n_136, n_134, n_132}));
  fx68k_mux_1834 mux_ccrMask_780_16(.ctl ({n_127, col[1], n_129,
       n_130}), .in_0 ({1'b0, ccrMask1[3], 1'b1, ccrMask1[1:0]}), .in_1
       ({n_139, n_137, n_135, n_133, n_131}), .in_2 ({n_140, 4'b1111}),
       .in_3 ({1'b0, n_138, n_136, n_134, n_132}), .z (ccrMask));
  or g1 (n_91, row[13], row[14]);
  not g9 (n_4, col[2]);
  nand g10 (n_149, n_4, n_7, col[1]);
  not g11 (n_97, n_149);
  not g12 (n_7, col[0]);
  nor g21 (n_43, row[9], row[3]);
  not g22 (n_113, n_43);
  nor g23 (n_44, row[2], row[5], row[10], row[12]);
  not g24 (n_114, n_44);
  nor g25 (n_45, row[6], row[7], row[11]);
  not g26 (n_115, n_45);
  nor g27 (n_46, row[4], row[8], row[13], row[14]);
  not g28 (n_116, n_46);
  nor g36 (n_127, col[2], col[1]);
  nor g37 (n_129, n_4, col[0]);
  nor g39 (n_130, n_4, n_7);
endmodule

module fx68k_bmux_1840(ctl, in_0, in_1, z);
  input ctl;
  input [31:0] in_0, in_1;
  output [31:0] z;
  wire ctl;
  wire [31:0] in_0, in_1;
  wire [31:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[31]), .data1 (in_1[31]), .z
       (z[31]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[30]), .data1 (in_1[30]), .z
       (z[30]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[29]), .data1 (in_1[29]), .z
       (z[29]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[28]), .data1 (in_1[28]), .z
       (z[28]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[27]), .data1 (in_1[27]), .z
       (z[27]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[26]), .data1 (in_1[26]), .z
       (z[26]));
  CDN_bmux2 g7(.sel0 (ctl), .data0 (in_0[25]), .data1 (in_1[25]), .z
       (z[25]));
  CDN_bmux2 g8(.sel0 (ctl), .data0 (in_0[24]), .data1 (in_1[24]), .z
       (z[24]));
  CDN_bmux2 g9(.sel0 (ctl), .data0 (in_0[23]), .data1 (in_1[23]), .z
       (z[23]));
  CDN_bmux2 g10(.sel0 (ctl), .data0 (in_0[22]), .data1 (in_1[22]), .z
       (z[22]));
  CDN_bmux2 g11(.sel0 (ctl), .data0 (in_0[21]), .data1 (in_1[21]), .z
       (z[21]));
  CDN_bmux2 g12(.sel0 (ctl), .data0 (in_0[20]), .data1 (in_1[20]), .z
       (z[20]));
  CDN_bmux2 g13(.sel0 (ctl), .data0 (in_0[19]), .data1 (in_1[19]), .z
       (z[19]));
  CDN_bmux2 g14(.sel0 (ctl), .data0 (in_0[18]), .data1 (in_1[18]), .z
       (z[18]));
  CDN_bmux2 g15(.sel0 (ctl), .data0 (in_0[17]), .data1 (in_1[17]), .z
       (z[17]));
  CDN_bmux2 g16(.sel0 (ctl), .data0 (in_0[16]), .data1 (in_1[16]), .z
       (z[16]));
  CDN_bmux2 g17(.sel0 (ctl), .data0 (in_0[15]), .data1 (in_1[15]), .z
       (z[15]));
  CDN_bmux2 g18(.sel0 (ctl), .data0 (in_0[14]), .data1 (in_1[14]), .z
       (z[14]));
  CDN_bmux2 g19(.sel0 (ctl), .data0 (in_0[13]), .data1 (in_1[13]), .z
       (z[13]));
  CDN_bmux2 g20(.sel0 (ctl), .data0 (in_0[12]), .data1 (in_1[12]), .z
       (z[12]));
  CDN_bmux2 g21(.sel0 (ctl), .data0 (in_0[11]), .data1 (in_1[11]), .z
       (z[11]));
  CDN_bmux2 g22(.sel0 (ctl), .data0 (in_0[10]), .data1 (in_1[10]), .z
       (z[10]));
  CDN_bmux2 g23(.sel0 (ctl), .data0 (in_0[9]), .data1 (in_1[9]), .z
       (z[9]));
  CDN_bmux2 g24(.sel0 (ctl), .data0 (in_0[8]), .data1 (in_1[8]), .z
       (z[8]));
  CDN_bmux2 g25(.sel0 (ctl), .data0 (in_0[7]), .data1 (in_1[7]), .z
       (z[7]));
  CDN_bmux2 g26(.sel0 (ctl), .data0 (in_0[6]), .data1 (in_1[6]), .z
       (z[6]));
  CDN_bmux2 g27(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g28(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g29(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g30(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g31(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g32(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_aluShifter(data, isByte, isLong, swapWords, dir, cin,
     result);
  input [31:0] data;
  input isByte, isLong, swapWords, dir, cin;
  output [31:0] result;
  wire [31:0] data;
  wire isByte, isLong, swapWords, dir, cin;
  wire [31:0] result;
  wire [31:0] tdata;
  wire n_1, n_2, n_3, n_7, n_10, n_11, n_12, n_13;
  wire n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21;
  wire n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_76;
  fx68k_bmux_1503 mux_tdata_504_20(.ctl (n_3), .in_0 (data[16]), .in_1
       (cin), .z (n_7));
  fx68k_bmux_1520 mux_tdata_502_14(.ctl (n_2), .in_0 ({n_7, data[8]}),
       .in_1 ({data[16], cin}), .z ({tdata[16], tdata[8]}));
  fx68k_bmux_1840 mux_result_516_12(.ctl (dir), .in_0 ({data[30:17],
       tdata[16], data[15:9], tdata[8], data[7:0], cin}), .in_1 ({cin,
       data[31:17], tdata[16], data[15:9], tdata[8], data[7:1]}), .z
       ({n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32,
       n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22,
       n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12,
       n_11, n_10}));
  fx68k_bmux_1840 mux_result_513_12(.ctl (swapWords), .in_0 ({n_41,
       n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31,
       n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21,
       n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11,
       n_10}), .in_1 ({data[30:17], tdata[16], cin, data[14:9],
       tdata[8], data[7:0], data[31]}), .z ({n_73, n_72, n_71, n_70,
       n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60,
       n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50,
       n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42}));
  fx68k_bmux_1840 mux_result_511_17(.ctl (n_1), .in_0 ({n_73, n_72,
       n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62,
       n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, n_52,
       n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42}),
       .in_1 ({data[0], data[31:17], cin, data[15:9], tdata[8],
       data[7:1]}), .z (result));
  and g1 (n_2, isByte, dir);
  and g3 (n_3, n_76, dir);
  and g4 (n_1, swapWords, dir);
  not g10 (n_76, isLong);
endmodule

module fx68k_add_unsigned(A, B, Z);
  input [7:0] A;
  input [8:0] B;
  output [8:0] Z;
  wire [7:0] A;
  wire [8:0] B;
  wire [8:0] Z;
  wire n_28, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46;
  wire n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62;
  wire n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_84, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_28, A[0], B[0]);
  nor g6 (n_32, A[1], B[1]);
  nand g7 (n_35, A[1], B[1]);
  nor g8 (n_42, A[2], B[2]);
  nand g9 (n_37, A[2], B[2]);
  nor g10 (n_38, A[3], B[3]);
  nand g11 (n_39, A[3], B[3]);
  nor g12 (n_48, A[4], B[4]);
  nand g13 (n_43, A[4], B[4]);
  nor g14 (n_44, A[5], B[5]);
  nand g15 (n_45, A[5], B[5]);
  nor g16 (n_54, A[6], B[6]);
  nand g17 (n_49, A[6], B[6]);
  nor g18 (n_50, A[7], B[7]);
  nand g19 (n_51, A[7], B[7]);
  not g22 (n_34, n_32);
  nand g23 (n_36, n_33, n_34);
  nand g24 (n_55, n_35, n_36);
  nor g25 (n_40, n_37, n_38);
  not g26 (n_41, n_39);
  nor g27 (n_59, n_40, n_41);
  nor g28 (n_58, n_42, n_38);
  nor g29 (n_46, n_43, n_44);
  not g30 (n_47, n_45);
  nor g31 (n_61, n_46, n_47);
  nor g32 (n_64, n_48, n_44);
  nor g33 (n_52, n_49, n_50);
  not g34 (n_53, n_51);
  nor g35 (n_68, n_52, n_53);
  nor g36 (n_66, n_54, n_50);
  not g37 (n_56, n_42);
  nand g38 (n_57, n_55, n_56);
  nand g39 (n_91, n_37, n_57);
  nand g40 (n_60, n_58, n_55);
  nand g41 (n_71, n_59, n_60);
  nor g42 (n_62, n_54, n_61);
  not g43 (n_63, n_49);
  nor g44 (n_77, n_62, n_63);
  not g45 (n_65, n_54);
  nand g46 (n_75, n_64, n_65);
  not g47 (n_67, n_66);
  nor g48 (n_69, n_61, n_67);
  not g49 (n_70, n_68);
  nor g50 (n_81, n_69, n_70);
  nand g51 (n_79, n_64, n_66);
  not g52 (n_72, n_48);
  nand g53 (n_73, n_71, n_72);
  nand g54 (n_95, n_43, n_73);
  nand g55 (n_74, n_64, n_71);
  nand g56 (n_97, n_61, n_74);
  not g57 (n_76, n_75);
  nand g58 (n_78, n_71, n_76);
  nand g59 (n_100, n_77, n_78);
  not g60 (n_80, n_79);
  nand g61 (n_82, n_71, n_80);
  nand g62 (n_84, n_81, n_82);
  nand g66 (n_88, n_34, n_35);
  xnor g67 (Z[1], n_33, n_88);
  nand g68 (n_89, n_56, n_37);
  xnor g69 (Z[2], n_55, n_89);
  not g70 (n_90, n_38);
  nand g71 (n_92, n_90, n_39);
  xnor g72 (Z[3], n_91, n_92);
  nand g73 (n_93, n_72, n_43);
  xnor g74 (Z[4], n_71, n_93);
  not g75 (n_94, n_44);
  nand g76 (n_96, n_94, n_45);
  xnor g77 (Z[5], n_95, n_96);
  nand g78 (n_98, n_65, n_49);
  xnor g79 (Z[6], n_97, n_98);
  not g80 (n_99, n_50);
  nand g81 (n_101, n_99, n_51);
  xnor g82 (Z[7], n_100, n_101);
  xnor g84 (Z[8], n_84, n_102);
  not g87 (n_33, n_28);
  not g88 (n_102, B[8]);
endmodule

module fx68k_sub_unsigned(A, B, Z);
  input [7:0] A;
  input [8:0] B;
  output [8:0] Z;
  wire [7:0] A;
  wire [8:0] B;
  wire [8:0] Z;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_41, n_43, n_44, n_45, n_46, n_47, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_95, n_99, n_100, n_101;
  wire n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109;
  wire n_110, n_111, n_112, n_114;
  not g3 (n_31, B[7]);
  not g4 (n_32, B[6]);
  not g5 (n_33, B[5]);
  not g6 (n_34, B[4]);
  not g7 (n_35, B[3]);
  not g8 (n_36, B[2]);
  not g9 (n_37, B[1]);
  not g10 (n_38, B[0]);
  xor g12 (n_114, A[0], n_38);
  nand g15 (n_44, n_41, B[0]);
  nor g16 (n_43, A[1], n_37);
  nand g17 (n_46, A[1], n_37);
  nor g18 (n_53, A[2], n_36);
  nand g19 (n_48, A[2], n_36);
  nor g20 (n_49, A[3], n_35);
  nand g21 (n_50, A[3], n_35);
  nor g22 (n_59, A[4], n_34);
  nand g23 (n_54, A[4], n_34);
  nor g24 (n_55, A[5], n_33);
  nand g25 (n_56, A[5], n_33);
  nor g26 (n_65, A[6], n_32);
  nand g27 (n_60, A[6], n_32);
  nor g28 (n_61, A[7], n_31);
  nand g29 (n_62, A[7], n_31);
  not g32 (n_45, n_43);
  nand g33 (n_47, n_44, n_45);
  nand g34 (n_66, n_46, n_47);
  nor g35 (n_51, n_48, n_49);
  not g36 (n_52, n_50);
  nor g37 (n_70, n_51, n_52);
  nor g38 (n_69, n_53, n_49);
  nor g39 (n_57, n_54, n_55);
  not g40 (n_58, n_56);
  nor g41 (n_72, n_57, n_58);
  nor g42 (n_75, n_59, n_55);
  nor g43 (n_63, n_60, n_61);
  not g44 (n_64, n_62);
  nor g45 (n_79, n_63, n_64);
  nor g46 (n_77, n_65, n_61);
  not g47 (n_67, n_53);
  nand g48 (n_68, n_66, n_67);
  nand g49 (n_102, n_48, n_68);
  nand g50 (n_71, n_69, n_66);
  nand g51 (n_82, n_70, n_71);
  nor g52 (n_73, n_65, n_72);
  not g53 (n_74, n_60);
  nor g54 (n_88, n_73, n_74);
  not g55 (n_76, n_65);
  nand g56 (n_86, n_75, n_76);
  not g57 (n_78, n_77);
  nor g58 (n_80, n_72, n_78);
  not g59 (n_81, n_79);
  nor g60 (n_92, n_80, n_81);
  nand g61 (n_90, n_75, n_77);
  not g62 (n_83, n_59);
  nand g63 (n_84, n_82, n_83);
  nand g64 (n_106, n_54, n_84);
  nand g65 (n_85, n_75, n_82);
  nand g66 (n_108, n_72, n_85);
  not g67 (n_87, n_86);
  nand g68 (n_89, n_82, n_87);
  nand g69 (n_111, n_88, n_89);
  not g70 (n_91, n_90);
  nand g71 (n_93, n_82, n_91);
  nand g72 (n_95, n_92, n_93);
  nand g76 (n_99, n_45, n_46);
  xnor g77 (Z[1], n_44, n_99);
  nand g78 (n_100, n_67, n_48);
  xnor g79 (Z[2], n_66, n_100);
  not g80 (n_101, n_49);
  nand g81 (n_103, n_101, n_50);
  xnor g82 (Z[3], n_102, n_103);
  nand g83 (n_104, n_83, n_54);
  xnor g84 (Z[4], n_82, n_104);
  not g85 (n_105, n_55);
  nand g86 (n_107, n_105, n_56);
  xnor g87 (Z[5], n_106, n_107);
  nand g88 (n_109, n_76, n_60);
  xnor g89 (Z[6], n_108, n_109);
  not g90 (n_110, n_61);
  nand g91 (n_112, n_110, n_62);
  xnor g92 (Z[7], n_111, n_112);
  xnor g94 (Z[8], n_95, B[8]);
  not g96 (n_41, A[0]);
  not g97 (Z[0], n_114);
endmodule

module fx68k_add_unsigned_1844(A, B, Z);
  input [4:0] A, B;
  output [4:0] Z;
  wire [4:0] A, B;
  wire [4:0] Z;
  wire n_17, n_20, n_21, n_22, n_23, n_24, n_25, n_26;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_42, n_43;
  wire n_44, n_45, n_46, n_47;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_17, A[0], B[0]);
  nor g6 (n_20, A[1], B[1]);
  nand g7 (n_23, A[1], B[1]);
  nor g8 (n_30, A[2], B[2]);
  nand g9 (n_25, A[2], B[2]);
  nor g10 (n_26, A[3], B[3]);
  nand g11 (n_27, A[3], B[3]);
  nor g12 (n_37, A[4], B[4]);
  nand g13 (n_40, A[4], B[4]);
  not g14 (n_22, n_20);
  nand g15 (n_24, n_21, n_22);
  nand g16 (n_31, n_23, n_24);
  nor g17 (n_28, n_25, n_26);
  not g18 (n_29, n_27);
  nor g19 (n_35, n_28, n_29);
  nor g20 (n_34, n_30, n_26);
  not g21 (n_32, n_30);
  nand g22 (n_33, n_31, n_32);
  nand g23 (n_45, n_25, n_33);
  nand g24 (n_36, n_34, n_31);
  nand g25 (n_38, n_35, n_36);
  not g26 (n_39, n_37);
  nand g29 (n_42, n_22, n_23);
  xnor g30 (Z[1], n_21, n_42);
  nand g31 (n_43, n_32, n_25);
  xnor g32 (Z[2], n_31, n_43);
  not g33 (n_44, n_26);
  nand g34 (n_46, n_44, n_27);
  xnor g35 (Z[3], n_45, n_46);
  nand g36 (n_47, n_39, n_40);
  xnor g37 (Z[4], n_38, n_47);
  not g39 (n_21, n_17);
endmodule

module fx68k_sub_unsigned_1846(A, B, Z);
  input [4:0] A, B;
  output [4:0] Z;
  wire [4:0] A, B;
  wire [4:0] Z;
  wire n_18, n_19, n_20, n_21, n_22, n_25, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_49, n_50, n_51, n_52, n_53;
  wire n_54, n_55;
  not g2 (n_18, B[4]);
  not g3 (n_19, B[3]);
  not g4 (n_20, B[2]);
  not g5 (n_21, B[1]);
  not g6 (n_22, B[0]);
  xor g8 (n_55, A[0], n_22);
  nand g11 (n_28, n_25, B[0]);
  nor g12 (n_27, A[1], n_21);
  nand g13 (n_30, A[1], n_21);
  nor g14 (n_37, A[2], n_20);
  nand g15 (n_32, A[2], n_20);
  nor g16 (n_33, A[3], n_19);
  nand g17 (n_34, A[3], n_19);
  nor g18 (n_44, A[4], n_18);
  nand g19 (n_47, A[4], n_18);
  not g20 (n_29, n_27);
  nand g21 (n_31, n_28, n_29);
  nand g22 (n_38, n_30, n_31);
  nor g23 (n_35, n_32, n_33);
  not g24 (n_36, n_34);
  nor g25 (n_42, n_35, n_36);
  nor g26 (n_41, n_37, n_33);
  not g27 (n_39, n_37);
  nand g28 (n_40, n_38, n_39);
  nand g29 (n_52, n_32, n_40);
  nand g30 (n_43, n_41, n_38);
  nand g31 (n_45, n_42, n_43);
  not g32 (n_46, n_44);
  nand g35 (n_49, n_29, n_30);
  xnor g36 (Z[1], n_28, n_49);
  nand g37 (n_50, n_39, n_32);
  xnor g38 (Z[2], n_38, n_50);
  not g39 (n_51, n_33);
  nand g40 (n_53, n_51, n_34);
  xnor g41 (Z[3], n_52, n_53);
  nand g42 (n_54, n_46, n_47);
  xnor g43 (Z[4], n_45, n_54);
  not g45 (n_25, A[0]);
  not g46 (Z[0], n_55);
endmodule

module fx68k_bmux_1854(ctl, in_0, in_1, z);
  input ctl;
  input [4:0] in_0, in_1;
  output [4:0] z;
  wire ctl;
  wire [4:0] in_0, in_1;
  wire [4:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_bmux_1855(ctl, in_0, in_1, z);
  input ctl;
  input [8:0] in_0, in_1;
  output [8:0] z;
  wire ctl;
  wire [8:0] in_0, in_1;
  wire [8:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[8]), .data1 (in_1[8]), .z
       (z[8]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[7]), .data1 (in_1[7]), .z
       (z[7]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[6]), .data1 (in_1[6]), .z
       (z[6]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g7(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g8(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g9(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_aluCorf(binResult, bAdd, cin, hCarry, bcdResult, dC, ov);
  input [7:0] binResult;
  input bAdd, cin, hCarry;
  output [7:0] bcdResult;
  output dC, ov;
  wire [7:0] binResult;
  wire bAdd, cin, hCarry;
  wire [7:0] bcdResult;
  wire dC, ov;
  wire [4:0] hNib;
  wire [8:0] htemp;
  wire highC, lowC, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_85, n_87, n_89, n_90, n_91, n_97;
  wire n_98, n_100, n_102, n_103, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, \nib[1]_119 ,
       \nib[2]_120 ;
  wire \nib[3]_121 ;
  fx68k_add_unsigned add_467_31(.A (binResult), .B ({6'b000000, n_110,
       n_109, 1'b0}), .Z ({n_90, \nib[3]_121 , \nib[2]_120 ,
       \nib[1]_119 , n_82, n_80, n_78, n_76, n_74}));
  fx68k_sub_unsigned sub_472_31(.A (binResult), .B ({6'b000000, n_112,
       n_111, 1'b0}), .Z ({n_91, n_89, n_87, n_85, n_83, n_81, n_79,
       n_77, n_75}));
  fx68k_add_unsigned_1844 add_468_23(.A ({n_90, \nib[3]_121 ,
       \nib[2]_120 , \nib[1]_119 , n_82}), .B ({2'b00, n_114, n_113,
       1'b0}), .Z ({n_72, n_70, n_68, n_66, n_64}));
  fx68k_sub_unsigned_1846 sub_473_23(.A ({n_91, n_89, n_87, n_85,
       n_83}), .B ({2'b00, n_116, n_115, 1'b0}), .Z ({n_73, n_71, n_69,
       n_67, n_65}));
  fx68k_bmux_1503 mux_462_25(.ctl (bAdd), .in_0 (1'b0), .in_1 (n_60),
       .z (n_97));
  fx68k_bmux_1520 mux_467_34(.ctl (lowC), .in_0 (2'b00), .in_1 (2'b11),
       .z ({n_110, n_109}));
  fx68k_bmux_1503 mux_463_22(.ctl (bAdd), .in_0 (1'b0), .in_1 (n_61),
       .z (n_100));
  fx68k_bmux_1520 mux_468_26(.ctl (highC), .in_0 (2'b00), .in_1
       (2'b11), .z ({n_114, n_113}));
  fx68k_bmux_1520 mux_472_34(.ctl (lowC), .in_0 (2'b00), .in_1 (2'b11),
       .z ({n_112, n_111}));
  fx68k_bmux_1520 mux_473_26(.ctl (highC), .in_0 (2'b00), .in_1
       (2'b11), .z ({n_116, n_115}));
  fx68k_bmux_1503 mux_ov_466_7(.ctl (bAdd), .in_0 (n_63), .in_1 (n_62),
       .z (ov));
  fx68k_bmux_1854 mux_hNib_466_7(.ctl (bAdd), .in_0 ({n_73, n_71, n_69,
       n_67, n_65}), .in_1 ({n_72, n_70, n_68, n_66, n_64}), .z
       ({hNib[4], bcdResult[7:4]}));
  fx68k_bmux_1855 mux_htemp_466_7(.ctl (bAdd), .in_0 ({n_91, n_89,
       n_87, n_85, n_83, n_81, n_79, n_77, n_75}), .in_1 ({n_90,
       \nib[3]_121 , \nib[2]_120 , \nib[1]_119 , n_82, n_80, n_78,
       n_76, n_74}), .z ({htemp[8:4], bcdResult[3:0]}));
  or g1 (lowC, hCarry, n_97);
  or g2 (n_61, n_98, n_90);
  or g3 (highC, cin, n_100);
  not g4 (n_102, binResult[7]);
  and g5 (n_62, n_70, n_102);
  not g6 (n_103, n_71);
  and g7 (n_63, n_103, binResult[7]);
  or g8 (dC, hNib[4], cin);
  or g12 (n_117, binResult[2], binResult[1]);
  and g13 (n_60, binResult[3], n_117);
  or g14 (n_118, \nib[2]_120 , \nib[1]_119 );
  and g15 (n_98, \nib[3]_121 , n_118);
endmodule

module fx68k_and_op(A, B, Z);
  input [15:0] A, B;
  output [15:0] Z;
  wire [15:0] A, B;
  wire [15:0] Z;
  and g1 (Z[0], A[0], B[0]);
  and g2 (Z[1], A[1], B[1]);
  and g3 (Z[2], A[2], B[2]);
  and g4 (Z[3], A[3], B[3]);
  and g5 (Z[4], A[4], B[4]);
  and g6 (Z[5], A[5], B[5]);
  and g7 (Z[6], A[6], B[6]);
  and g8 (Z[7], A[7], B[7]);
  and g9 (Z[8], A[8], B[8]);
  and g10 (Z[9], A[9], B[9]);
  and g11 (Z[10], A[10], B[10]);
  and g12 (Z[11], A[11], B[11]);
  and g13 (Z[12], A[12], B[12]);
  and g14 (Z[13], A[13], B[13]);
  and g15 (Z[14], A[14], B[14]);
  and g16 (Z[15], A[15], B[15]);
endmodule

module fx68k_or_op_1132(A, B, Z);
  input [15:0] A, B;
  output [15:0] Z;
  wire [15:0] A, B;
  wire [15:0] Z;
  or g1 (Z[0], A[0], B[0]);
  or g2 (Z[1], A[1], B[1]);
  or g3 (Z[2], A[2], B[2]);
  or g4 (Z[3], A[3], B[3]);
  or g5 (Z[4], A[4], B[4]);
  or g6 (Z[5], A[5], B[5]);
  or g7 (Z[6], A[6], B[6]);
  or g8 (Z[7], A[7], B[7]);
  or g9 (Z[8], A[8], B[8]);
  or g10 (Z[9], A[9], B[9]);
  or g11 (Z[10], A[10], B[10]);
  or g12 (Z[11], A[11], B[11]);
  or g13 (Z[12], A[12], B[12]);
  or g14 (Z[13], A[13], B[13]);
  or g15 (Z[14], A[14], B[14]);
  or g16 (Z[15], A[15], B[15]);
endmodule

module fx68k_xor_op(A, B, Z);
  input [15:0] A, B;
  output [15:0] Z;
  wire [15:0] A, B;
  wire [15:0] Z;
  xor g1 (Z[0], A[0], B[0]);
  xor g2 (Z[1], A[1], B[1]);
  xor g3 (Z[2], A[2], B[2]);
  xor g4 (Z[3], A[3], B[3]);
  xor g5 (Z[4], A[4], B[4]);
  xor g6 (Z[5], A[5], B[5]);
  xor g7 (Z[6], A[6], B[6]);
  xor g8 (Z[7], A[7], B[7]);
  xor g9 (Z[8], A[8], B[8]);
  xor g10 (Z[9], A[9], B[9]);
  xor g11 (Z[10], A[10], B[10]);
  xor g12 (Z[11], A[11], B[11]);
  xor g13 (Z[12], A[12], B[12]);
  xor g14 (Z[13], A[13], B[13]);
  xor g15 (Z[14], A[14], B[14]);
  xor g16 (Z[15], A[15], B[15]);
endmodule

module fx68k_or_op_1133(A, Z);
  input [7:0] A;
  output Z;
  wire [7:0] A;
  wire Z;
  wire n_9, n_10;
  nor g1 (n_10, A[7], A[6], A[5], A[4]);
  nor g2 (n_9, A[3], A[2], A[1], A[0]);
  nand g3 (Z, n_9, n_10);
endmodule

module fx68k_or_op_1134(A, Z);
  input [15:0] A;
  output Z;
  wire [15:0] A;
  wire Z;
  wire n_17, n_18, n_19, n_20;
  nor g1 (n_17, A[15], A[14], A[13], A[12]);
  nor g2 (n_18, A[11], A[10], A[9], A[8]);
  nor g3 (n_19, A[7], A[6], A[5], A[4]);
  nor g4 (n_20, A[3], A[2], A[1], A[0]);
  nand g5 (Z, n_17, n_18, n_19, n_20);
endmodule

module fx68k_and_op_1135(A, B, Z);
  input [4:0] A, B;
  output [4:0] Z;
  wire [4:0] A, B;
  wire [4:0] Z;
  and g1 (Z[0], A[0], B[0]);
  and g2 (Z[1], A[1], B[1]);
  and g3 (Z[2], A[2], B[2]);
  and g4 (Z[3], A[3], B[3]);
  and g5 (Z[4], A[4], B[4]);
endmodule

module fx68k_not_op(A, Z);
  input [4:0] A;
  output [4:0] Z;
  wire [4:0] A;
  wire [4:0] Z;
  not g1 (Z[4], A[4]);
  not g2 (Z[3], A[3]);
  not g3 (Z[2], A[2]);
  not g4 (Z[1], A[1]);
  not g5 (Z[0], A[0]);
endmodule

module fx68k_and_op_1136(A, B, Z);
  input [4:0] A, B;
  output [4:0] Z;
  wire [4:0] A, B;
  wire [4:0] Z;
  and g1 (Z[0], A[0], B[0]);
  and g2 (Z[1], A[1], B[1]);
  and g3 (Z[2], A[2], B[2]);
  and g4 (Z[3], A[3], B[3]);
  and g5 (Z[4], A[4], B[4]);
endmodule

module fx68k_or_op_1137(A, B, Z);
  input [4:0] A, B;
  output [4:0] Z;
  wire [4:0] A, B;
  wire [4:0] Z;
  or g1 (Z[0], A[0], B[0]);
  or g2 (Z[1], A[1], B[1]);
  or g3 (Z[2], A[2], B[2]);
  or g4 (Z[3], A[3], B[3]);
  or g5 (Z[4], A[4], B[4]);
endmodule

module fx68k_or_op_1138(A, Z);
  input [2:0] A;
  output Z;
  wire [2:0] A;
  wire Z;
  wire n_4;
  nor g1 (n_4, A[2], A[1], A[0]);
  not g2 (Z, n_4);
endmodule

module fx68k_add_unsigned_1865(A, B, Z);
  input [8:0] A, B;
  output [9:0] Z;
  wire [8:0] A, B;
  wire [9:0] Z;
  wire n_30, n_33, n_34, n_35, n_36, n_37, n_38, n_39;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_30, A[0], B[0]);
  nor g6 (n_33, A[1], B[1]);
  nand g7 (n_36, A[1], B[1]);
  nor g8 (n_43, A[2], B[2]);
  nand g9 (n_38, A[2], B[2]);
  nor g10 (n_39, A[3], B[3]);
  nand g11 (n_40, A[3], B[3]);
  nor g12 (n_49, A[4], B[4]);
  nand g13 (n_44, A[4], B[4]);
  nor g14 (n_45, A[5], B[5]);
  nand g15 (n_46, A[5], B[5]);
  nor g16 (n_55, A[6], B[6]);
  nand g17 (n_50, A[6], B[6]);
  nor g18 (n_51, A[7], B[7]);
  nand g19 (n_52, A[7], B[7]);
  nor g20 (n_84, A[8], B[8]);
  nand g21 (n_87, A[8], B[8]);
  not g22 (n_35, n_33);
  nand g23 (n_37, n_34, n_35);
  nand g24 (n_56, n_36, n_37);
  nor g25 (n_41, n_38, n_39);
  not g26 (n_42, n_40);
  nor g27 (n_60, n_41, n_42);
  nor g28 (n_59, n_43, n_39);
  nor g29 (n_47, n_44, n_45);
  not g30 (n_48, n_46);
  nor g31 (n_62, n_47, n_48);
  nor g32 (n_65, n_49, n_45);
  nor g33 (n_53, n_50, n_51);
  not g34 (n_54, n_52);
  nor g35 (n_69, n_53, n_54);
  nor g36 (n_67, n_55, n_51);
  not g37 (n_57, n_43);
  nand g38 (n_58, n_56, n_57);
  nand g39 (n_92, n_38, n_58);
  nand g40 (n_61, n_59, n_56);
  nand g41 (n_72, n_60, n_61);
  nor g42 (n_63, n_55, n_62);
  not g43 (n_64, n_50);
  nor g44 (n_78, n_63, n_64);
  not g45 (n_66, n_55);
  nand g46 (n_76, n_65, n_66);
  not g47 (n_68, n_67);
  nor g48 (n_70, n_62, n_68);
  not g49 (n_71, n_69);
  nor g50 (n_82, n_70, n_71);
  nand g51 (n_80, n_65, n_67);
  not g52 (n_73, n_49);
  nand g53 (n_74, n_72, n_73);
  nand g54 (n_96, n_44, n_74);
  nand g55 (n_75, n_65, n_72);
  nand g56 (n_98, n_62, n_75);
  not g57 (n_77, n_76);
  nand g58 (n_79, n_72, n_77);
  nand g59 (n_101, n_78, n_79);
  not g60 (n_81, n_80);
  nand g61 (n_83, n_72, n_81);
  nand g62 (n_85, n_82, n_83);
  not g63 (n_86, n_84);
  nand g64 (n_88, n_85, n_86);
  nand g65 (Z[9], n_87, n_88);
  nand g66 (n_89, n_35, n_36);
  xnor g67 (Z[1], n_34, n_89);
  nand g68 (n_90, n_57, n_38);
  xnor g69 (Z[2], n_56, n_90);
  not g70 (n_91, n_39);
  nand g71 (n_93, n_91, n_40);
  xnor g72 (Z[3], n_92, n_93);
  nand g73 (n_94, n_73, n_44);
  xnor g74 (Z[4], n_72, n_94);
  not g75 (n_95, n_45);
  nand g76 (n_97, n_95, n_46);
  xnor g77 (Z[5], n_96, n_97);
  nand g78 (n_99, n_66, n_50);
  xnor g79 (Z[6], n_98, n_99);
  not g80 (n_100, n_51);
  nand g81 (n_102, n_100, n_52);
  xnor g82 (Z[7], n_101, n_102);
  nand g83 (n_103, n_86, n_87);
  xnor g84 (Z[8], n_85, n_103);
  not g86 (n_34, n_30);
endmodule

module fx68k_add_unsigned_1867(A, B, Z);
  input [9:0] A;
  input B;
  output [10:0] Z;
  wire [9:0] A;
  wire B;
  wire [10:0] Z;
  wire n_24, n_37, n_40, n_42, n_46, n_48, n_52, n_54;
  wire n_58, n_60, n_64, n_65, n_67, n_68, n_70, n_74;
  wire n_76, n_81, n_83, n_84, n_85, n_86, n_88, n_89;
  wire n_90, n_92, n_93, n_95, n_96, n_98, n_99, n_102;
  wire n_106, n_108, n_111, n_115;
  xor g1 (Z[0], A[0], B);
  nand g2 (n_24, A[0], B);
  nand g25 (n_40, n_37, A[1]);
  nor g30 (n_68, n_46, n_42);
  nor g34 (n_74, n_52, n_48);
  nor g38 (n_76, n_58, n_54);
  nor g42 (n_96, n_64, n_60);
  nand g44 (n_67, n_65, A[2]);
  nand g46 (n_70, n_68, n_65);
  nand g52 (n_85, n_74, A[6]);
  nand g57 (n_89, n_74, n_76);
  nand g59 (n_83, n_81, A[4]);
  nand g61 (n_84, n_74, n_81);
  not g63 (n_86, n_85);
  nand g64 (n_88, n_81, n_86);
  not g66 (n_90, n_89);
  nand g67 (n_92, n_81, n_90);
  nand g70 (n_95, n_93, A[8]);
  nand g72 (n_98, n_96, n_93);
  xnor g75 (Z[1], n_37, n_99);
  xnor g77 (Z[2], n_65, n_46);
  xnor g80 (Z[3], n_102, n_42);
  xnor g82 (Z[4], n_81, n_52);
  xnor g85 (Z[5], n_106, n_48);
  xnor g87 (Z[6], n_108, n_58);
  xnor g90 (Z[7], n_111, n_54);
  xnor g92 (Z[8], n_93, n_64);
  xnor g95 (Z[9], n_115, n_60);
  not g98 (n_46, A[2]);
  not g99 (n_42, A[3]);
  not g100 (n_52, A[4]);
  not g101 (n_48, A[5]);
  not g102 (n_58, A[6]);
  not g103 (n_54, A[7]);
  not g104 (n_64, A[8]);
  not g105 (n_60, A[9]);
  not g106 (n_37, n_24);
  not g107 (n_99, A[1]);
  not g108 (n_65, n_40);
  not g109 (n_102, n_67);
  not g110 (n_81, n_70);
  not g111 (n_106, n_83);
  not g112 (n_108, n_84);
  not g113 (n_111, n_88);
  not g114 (n_93, n_92);
  not g115 (n_115, n_95);
  not g116 (Z[10], n_98);
endmodule

module fx68k_sub_unsigned_1869(A, B, Z);
  input [8:0] A, B;
  output [9:0] Z;
  wire [8:0] A, B;
  wire [9:0] Z;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_39, n_40, n_41, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114;
  not g2 (n_31, B[8]);
  not g3 (n_32, B[7]);
  not g4 (n_33, B[6]);
  not g5 (n_34, B[5]);
  not g6 (n_35, B[4]);
  not g7 (n_36, B[3]);
  not g8 (n_37, B[2]);
  not g9 (n_38, B[1]);
  not g10 (n_39, B[0]);
  not g11 (Z[9], n_40);
  xor g12 (n_114, A[0], n_39);
  nand g15 (n_44, n_41, B[0]);
  nor g16 (n_43, A[1], n_38);
  nand g17 (n_46, A[1], n_38);
  nor g18 (n_53, A[2], n_37);
  nand g19 (n_48, A[2], n_37);
  nor g20 (n_49, A[3], n_36);
  nand g21 (n_50, A[3], n_36);
  nor g22 (n_59, A[4], n_35);
  nand g23 (n_54, A[4], n_35);
  nor g24 (n_55, A[5], n_34);
  nand g25 (n_56, A[5], n_34);
  nor g26 (n_65, A[6], n_33);
  nand g27 (n_60, A[6], n_33);
  nor g28 (n_61, A[7], n_32);
  nand g29 (n_62, A[7], n_32);
  nor g30 (n_94, A[8], n_31);
  nand g31 (n_97, A[8], n_31);
  not g32 (n_45, n_43);
  nand g33 (n_47, n_44, n_45);
  nand g34 (n_66, n_46, n_47);
  nor g35 (n_51, n_48, n_49);
  not g36 (n_52, n_50);
  nor g37 (n_70, n_51, n_52);
  nor g38 (n_69, n_53, n_49);
  nor g39 (n_57, n_54, n_55);
  not g40 (n_58, n_56);
  nor g41 (n_72, n_57, n_58);
  nor g42 (n_75, n_59, n_55);
  nor g43 (n_63, n_60, n_61);
  not g44 (n_64, n_62);
  nor g45 (n_79, n_63, n_64);
  nor g46 (n_77, n_65, n_61);
  not g47 (n_67, n_53);
  nand g48 (n_68, n_66, n_67);
  nand g49 (n_102, n_48, n_68);
  nand g50 (n_71, n_69, n_66);
  nand g51 (n_82, n_70, n_71);
  nor g52 (n_73, n_65, n_72);
  not g53 (n_74, n_60);
  nor g54 (n_88, n_73, n_74);
  not g55 (n_76, n_65);
  nand g56 (n_86, n_75, n_76);
  not g57 (n_78, n_77);
  nor g58 (n_80, n_72, n_78);
  not g59 (n_81, n_79);
  nor g60 (n_92, n_80, n_81);
  nand g61 (n_90, n_75, n_77);
  not g62 (n_83, n_59);
  nand g63 (n_84, n_82, n_83);
  nand g64 (n_106, n_54, n_84);
  nand g65 (n_85, n_75, n_82);
  nand g66 (n_108, n_72, n_85);
  not g67 (n_87, n_86);
  nand g68 (n_89, n_82, n_87);
  nand g69 (n_111, n_88, n_89);
  not g70 (n_91, n_90);
  nand g71 (n_93, n_82, n_91);
  nand g72 (n_95, n_92, n_93);
  not g73 (n_96, n_94);
  nand g74 (n_98, n_95, n_96);
  nand g75 (n_40, n_97, n_98);
  nand g76 (n_99, n_45, n_46);
  xnor g77 (Z[1], n_44, n_99);
  nand g78 (n_100, n_67, n_48);
  xnor g79 (Z[2], n_66, n_100);
  not g80 (n_101, n_49);
  nand g81 (n_103, n_101, n_50);
  xnor g82 (Z[3], n_102, n_103);
  nand g83 (n_104, n_83, n_54);
  xnor g84 (Z[4], n_82, n_104);
  not g85 (n_105, n_55);
  nand g86 (n_107, n_105, n_56);
  xnor g87 (Z[5], n_106, n_107);
  nand g88 (n_109, n_76, n_60);
  xnor g89 (Z[6], n_108, n_109);
  not g90 (n_110, n_61);
  nand g91 (n_112, n_110, n_62);
  xnor g92 (Z[7], n_111, n_112);
  nand g93 (n_113, n_96, n_97);
  xnor g94 (Z[8], n_95, n_113);
  not g96 (n_41, A[0]);
  not g97 (Z[0], n_114);
endmodule

module fx68k_sub_signed(A, B, Z);
  input [9:0] A;
  input [1:0] B;
  output [16:0] Z;
  wire [9:0] A;
  wire [1:0] B;
  wire [16:0] Z;
  wire n_26, n_27, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_47, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  assign Z[10] = Z[16];
  assign Z[11] = Z[16];
  assign Z[12] = Z[16];
  assign Z[13] = Z[16];
  assign Z[14] = Z[16];
  assign Z[15] = Z[16];
  not g2 (n_26, B[0]);
  not g3 (n_27, B[1]);
  not g11 (n_35, A[9]);
  not g12 (Z[16], n_43);
  xor g13 (n_120, A[0], n_26);
  nand g16 (n_48, n_45, B[0]);
  nor g17 (n_47, A[1], n_27);
  nand g18 (n_50, A[1], n_27);
  nor g19 (n_57, A[2], n_27);
  nand g20 (n_52, A[2], n_27);
  nor g21 (n_53, A[3], n_27);
  nand g22 (n_54, A[3], n_27);
  nor g23 (n_40, A[4], n_27);
  nand g24 (n_58, A[4], n_27);
  nor g25 (n_36, A[5], n_27);
  nand g26 (n_37, A[5], n_27);
  nor g27 (n_61, A[6], n_27);
  nand g28 (n_41, A[6], n_27);
  nor g29 (n_42, A[7], n_27);
  nand g30 (n_59, A[7], n_27);
  nor g31 (n_67, A[8], n_27);
  nand g32 (n_62, A[8], n_27);
  nor g33 (n_63, n_35, B[1]);
  nand g34 (n_64, n_35, B[1]);
  not g35 (n_49, n_47);
  nand g36 (n_51, n_48, n_49);
  nand g37 (n_68, n_50, n_51);
  nor g38 (n_55, n_52, n_53);
  not g39 (n_56, n_54);
  nor g40 (n_72, n_55, n_56);
  nor g41 (n_71, n_57, n_53);
  nor g42 (n_38, n_58, n_36);
  not g43 (n_39, n_37);
  nor g44 (n_74, n_38, n_39);
  nor g45 (n_77, n_40, n_36);
  nor g46 (n_44, n_41, n_42);
  not g47 (n_60, n_59);
  nor g48 (n_81, n_44, n_60);
  nor g49 (n_79, n_61, n_42);
  nor g50 (n_65, n_62, n_63);
  not g51 (n_66, n_64);
  nor g52 (n_100, n_65, n_66);
  nor g53 (n_99, n_67, n_63);
  not g54 (n_69, n_57);
  nand g55 (n_70, n_68, n_69);
  nand g56 (n_105, n_52, n_70);
  nand g57 (n_73, n_71, n_68);
  nand g58 (n_84, n_72, n_73);
  nor g59 (n_75, n_61, n_74);
  not g60 (n_76, n_41);
  nor g61 (n_90, n_75, n_76);
  not g62 (n_78, n_61);
  nand g63 (n_88, n_77, n_78);
  not g64 (n_80, n_79);
  nor g65 (n_82, n_74, n_80);
  not g66 (n_83, n_81);
  nor g67 (n_94, n_82, n_83);
  nand g68 (n_92, n_77, n_79);
  not g69 (n_85, n_40);
  nand g70 (n_86, n_84, n_85);
  nand g71 (n_109, n_58, n_86);
  nand g72 (n_87, n_77, n_84);
  nand g73 (n_111, n_74, n_87);
  not g74 (n_89, n_88);
  nand g75 (n_91, n_84, n_89);
  nand g76 (n_114, n_90, n_91);
  not g77 (n_93, n_92);
  nand g78 (n_95, n_84, n_93);
  nand g79 (n_96, n_94, n_95);
  not g80 (n_97, n_67);
  nand g81 (n_98, n_96, n_97);
  nand g82 (n_118, n_62, n_98);
  nand g83 (n_101, n_99, n_96);
  nand g84 (n_43, n_100, n_101);
  nand g85 (n_102, n_49, n_50);
  xnor g86 (Z[1], n_48, n_102);
  nand g87 (n_103, n_69, n_52);
  xnor g88 (Z[2], n_68, n_103);
  not g89 (n_104, n_53);
  nand g90 (n_106, n_104, n_54);
  xnor g91 (Z[3], n_105, n_106);
  nand g92 (n_107, n_85, n_58);
  xnor g93 (Z[4], n_84, n_107);
  not g94 (n_108, n_36);
  nand g95 (n_110, n_108, n_37);
  xnor g96 (Z[5], n_109, n_110);
  nand g97 (n_112, n_78, n_41);
  xnor g98 (Z[6], n_111, n_112);
  not g99 (n_113, n_42);
  nand g100 (n_115, n_113, n_59);
  xnor g101 (Z[7], n_114, n_115);
  nand g102 (n_116, n_97, n_62);
  xnor g103 (Z[8], n_96, n_116);
  not g104 (n_117, n_63);
  nand g105 (n_119, n_117, n_64);
  xnor g106 (Z[9], n_118, n_119);
  not g108 (n_45, A[0]);
  not g109 (Z[0], n_120);
endmodule

module fx68k_add_unsigned_1871(A, B, Z);
  input [15:0] A, B;
  output [16:0] Z;
  wire [15:0] A, B;
  wire [16:0] Z;
  wire n_51, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_51, A[0], B[0]);
  nor g6 (n_54, A[1], B[1]);
  nand g7 (n_57, A[1], B[1]);
  nor g8 (n_64, A[2], B[2]);
  nand g9 (n_59, A[2], B[2]);
  nor g10 (n_60, A[3], B[3]);
  nand g11 (n_61, A[3], B[3]);
  nor g12 (n_70, A[4], B[4]);
  nand g13 (n_65, A[4], B[4]);
  nor g14 (n_66, A[5], B[5]);
  nand g15 (n_67, A[5], B[5]);
  nor g16 (n_76, A[6], B[6]);
  nand g17 (n_71, A[6], B[6]);
  nor g18 (n_72, A[7], B[7]);
  nand g19 (n_73, A[7], B[7]);
  nor g20 (n_82, A[8], B[8]);
  nand g21 (n_77, A[8], B[8]);
  nor g22 (n_78, A[9], B[9]);
  nand g23 (n_79, A[9], B[9]);
  nor g24 (n_88, A[10], B[10]);
  nand g25 (n_83, A[10], B[10]);
  nor g26 (n_84, A[11], B[11]);
  nand g27 (n_85, A[11], B[11]);
  nor g28 (n_94, A[12], B[12]);
  nand g29 (n_89, A[12], B[12]);
  nor g30 (n_90, A[13], B[13]);
  nand g31 (n_91, A[13], B[13]);
  nor g32 (n_100, A[14], B[14]);
  nand g33 (n_95, A[14], B[14]);
  nor g34 (n_96, A[15], B[15]);
  nand g35 (n_97, A[15], B[15]);
  not g36 (n_56, n_54);
  nand g37 (n_58, n_55, n_56);
  nand g38 (n_101, n_57, n_58);
  nor g39 (n_62, n_59, n_60);
  not g40 (n_63, n_61);
  nor g41 (n_105, n_62, n_63);
  nor g42 (n_104, n_64, n_60);
  nor g43 (n_68, n_65, n_66);
  not g44 (n_69, n_67);
  nor g45 (n_107, n_68, n_69);
  nor g46 (n_110, n_70, n_66);
  nor g47 (n_74, n_71, n_72);
  not g48 (n_75, n_73);
  nor g49 (n_114, n_74, n_75);
  nor g50 (n_112, n_76, n_72);
  nor g51 (n_80, n_77, n_78);
  not g52 (n_81, n_79);
  nor g53 (n_117, n_80, n_81);
  nor g54 (n_120, n_82, n_78);
  nor g55 (n_86, n_83, n_84);
  not g56 (n_87, n_85);
  nor g57 (n_124, n_86, n_87);
  nor g58 (n_122, n_88, n_84);
  nor g59 (n_92, n_89, n_90);
  not g60 (n_93, n_91);
  nor g61 (n_127, n_92, n_93);
  nor g62 (n_130, n_94, n_90);
  nor g63 (n_98, n_95, n_96);
  not g64 (n_99, n_97);
  nor g65 (n_134, n_98, n_99);
  nor g66 (n_132, n_100, n_96);
  not g67 (n_102, n_64);
  nand g68 (n_103, n_101, n_102);
  nand g69 (n_189, n_59, n_103);
  nand g70 (n_106, n_104, n_101);
  nand g71 (n_137, n_105, n_106);
  nor g72 (n_108, n_76, n_107);
  not g73 (n_109, n_71);
  nor g74 (n_143, n_108, n_109);
  not g75 (n_111, n_76);
  nand g76 (n_141, n_110, n_111);
  not g77 (n_113, n_112);
  nor g78 (n_115, n_107, n_113);
  not g79 (n_116, n_114);
  nor g80 (n_147, n_115, n_116);
  nand g81 (n_145, n_110, n_112);
  nor g82 (n_118, n_88, n_117);
  not g83 (n_119, n_83);
  nor g84 (n_170, n_118, n_119);
  not g85 (n_121, n_88);
  nand g86 (n_168, n_120, n_121);
  not g87 (n_123, n_122);
  nor g88 (n_125, n_117, n_123);
  not g89 (n_126, n_124);
  nor g90 (n_149, n_125, n_126);
  nand g91 (n_152, n_120, n_122);
  nor g92 (n_128, n_100, n_127);
  not g93 (n_129, n_95);
  nor g94 (n_157, n_128, n_129);
  not g95 (n_131, n_100);
  nand g96 (n_156, n_130, n_131);
  not g97 (n_133, n_132);
  nor g98 (n_135, n_127, n_133);
  not g99 (n_136, n_134);
  nor g100 (n_161, n_135, n_136);
  nand g101 (n_160, n_130, n_132);
  not g102 (n_138, n_70);
  nand g103 (n_139, n_137, n_138);
  nand g104 (n_193, n_65, n_139);
  nand g105 (n_140, n_110, n_137);
  nand g106 (n_195, n_107, n_140);
  not g107 (n_142, n_141);
  nand g108 (n_144, n_137, n_142);
  nand g109 (n_198, n_143, n_144);
  not g110 (n_146, n_145);
  nand g111 (n_148, n_137, n_146);
  nand g112 (n_164, n_147, n_148);
  nor g113 (n_150, n_94, n_149);
  not g114 (n_151, n_89);
  nor g115 (n_175, n_150, n_151);
  nor g116 (n_174, n_94, n_152);
  not g117 (n_153, n_130);
  nor g118 (n_154, n_149, n_153);
  not g119 (n_155, n_127);
  nor g120 (n_178, n_154, n_155);
  nor g121 (n_177, n_152, n_153);
  nor g122 (n_158, n_156, n_149);
  not g123 (n_159, n_157);
  nor g124 (n_181, n_158, n_159);
  nor g125 (n_180, n_152, n_156);
  nor g126 (n_162, n_160, n_149);
  not g127 (n_163, n_161);
  nor g128 (n_184, n_162, n_163);
  nor g129 (n_183, n_152, n_160);
  not g130 (n_165, n_82);
  nand g131 (n_166, n_164, n_165);
  nand g132 (n_202, n_77, n_166);
  nand g133 (n_167, n_120, n_164);
  nand g134 (n_204, n_117, n_167);
  not g135 (n_169, n_168);
  nand g136 (n_171, n_164, n_169);
  nand g137 (n_207, n_170, n_171);
  not g138 (n_172, n_152);
  nand g139 (n_173, n_164, n_172);
  nand g140 (n_210, n_149, n_173);
  nand g141 (n_176, n_174, n_164);
  nand g142 (n_213, n_175, n_176);
  nand g143 (n_179, n_177, n_164);
  nand g144 (n_215, n_178, n_179);
  nand g145 (n_182, n_180, n_164);
  nand g146 (n_218, n_181, n_182);
  nand g147 (n_185, n_183, n_164);
  nand g148 (Z[16], n_184, n_185);
  nand g149 (n_186, n_56, n_57);
  xnor g150 (Z[1], n_55, n_186);
  nand g151 (n_187, n_102, n_59);
  xnor g152 (Z[2], n_101, n_187);
  not g153 (n_188, n_60);
  nand g154 (n_190, n_188, n_61);
  xnor g155 (Z[3], n_189, n_190);
  nand g156 (n_191, n_138, n_65);
  xnor g157 (Z[4], n_137, n_191);
  not g158 (n_192, n_66);
  nand g159 (n_194, n_192, n_67);
  xnor g160 (Z[5], n_193, n_194);
  nand g161 (n_196, n_111, n_71);
  xnor g162 (Z[6], n_195, n_196);
  not g163 (n_197, n_72);
  nand g164 (n_199, n_197, n_73);
  xnor g165 (Z[7], n_198, n_199);
  nand g166 (n_200, n_165, n_77);
  xnor g167 (Z[8], n_164, n_200);
  not g168 (n_201, n_78);
  nand g169 (n_203, n_201, n_79);
  xnor g170 (Z[9], n_202, n_203);
  nand g171 (n_205, n_121, n_83);
  xnor g172 (Z[10], n_204, n_205);
  not g173 (n_206, n_84);
  nand g174 (n_208, n_206, n_85);
  xnor g175 (Z[11], n_207, n_208);
  not g176 (n_209, n_94);
  nand g177 (n_211, n_209, n_89);
  xnor g178 (Z[12], n_210, n_211);
  not g179 (n_212, n_90);
  nand g180 (n_214, n_212, n_91);
  xnor g181 (Z[13], n_213, n_214);
  nand g182 (n_216, n_131, n_95);
  xnor g183 (Z[14], n_215, n_216);
  not g184 (n_217, n_96);
  nand g185 (n_219, n_217, n_97);
  xnor g186 (Z[15], n_218, n_219);
  not g188 (n_55, n_51);
endmodule

module fx68k_add_unsigned_1873(A, B, Z);
  input [16:0] A;
  input B;
  output [16:0] Z;
  wire [16:0] A;
  wire B;
  wire [16:0] Z;
  wire n_37, n_57, n_60, n_62, n_66, n_68, n_72, n_74;
  wire n_78, n_80, n_84, n_86, n_90, n_92, n_96, n_98;
  wire n_102, n_103, n_105, n_106, n_108, n_112, n_114, n_122;
  wire n_124, n_132, n_134, n_139, n_141, n_142, n_143, n_144;
  wire n_146, n_147, n_148, n_150, n_154, n_155, n_158, n_162;
  wire n_166, n_168, n_169, n_170, n_171, n_173, n_174, n_175;
  wire n_176, n_178, n_179, n_181, n_182, n_184, n_185, n_187;
  wire n_189, n_193, n_196, n_200, n_202, n_205, n_209, n_211;
  wire n_214, n_217, n_220, n_222, n_225, n_227;
  xor g1 (Z[0], A[0], B);
  nand g2 (n_37, A[0], B);
  nand g39 (n_60, n_57, A[1]);
  nor g44 (n_106, n_66, n_62);
  nor g48 (n_112, n_72, n_68);
  nor g52 (n_114, n_78, n_74);
  nor g56 (n_122, n_84, n_80);
  nor g60 (n_124, n_90, n_86);
  nor g64 (n_132, n_96, n_92);
  nor g68 (n_134, n_102, n_98);
  nand g70 (n_105, n_103, A[2]);
  nand g72 (n_108, n_106, n_103);
  nand g78 (n_143, n_112, A[6]);
  nand g83 (n_147, n_112, n_114);
  nand g88 (n_170, n_122, A[10]);
  nand g93 (n_154, n_122, n_124);
  nand g98 (n_158, n_132, A[14]);
  nand g103 (n_162, n_132, n_134);
  nand g105 (n_141, n_139, A[4]);
  nand g107 (n_142, n_112, n_139);
  not g109 (n_144, n_143);
  nand g110 (n_146, n_139, n_144);
  not g112 (n_148, n_147);
  nand g113 (n_150, n_139, n_148);
  nor g118 (n_176, n_96, n_154);
  not g119 (n_155, n_132);
  nor g123 (n_179, n_154, n_155);
  nor g127 (n_182, n_154, n_158);
  nor g131 (n_185, n_154, n_162);
  nand g133 (n_168, n_166, A[8]);
  nand g135 (n_169, n_122, n_166);
  not g137 (n_171, n_170);
  nand g138 (n_173, n_166, n_171);
  not g140 (n_174, n_154);
  nand g141 (n_175, n_166, n_174);
  nand g143 (n_178, n_176, n_166);
  nand g145 (n_181, n_179, n_166);
  nand g147 (n_184, n_182, n_166);
  nand g149 (n_187, n_185, n_166);
  xnor g155 (Z[1], n_57, n_193);
  xnor g157 (Z[2], n_103, n_66);
  xnor g160 (Z[3], n_196, n_62);
  xnor g162 (Z[4], n_139, n_72);
  xnor g165 (Z[5], n_200, n_68);
  xnor g167 (Z[6], n_202, n_78);
  xnor g170 (Z[7], n_205, n_74);
  xnor g172 (Z[8], n_166, n_84);
  xnor g175 (Z[9], n_209, n_80);
  xnor g177 (Z[10], n_211, n_90);
  xnor g180 (Z[11], n_214, n_86);
  xnor g183 (Z[12], n_217, n_96);
  xnor g186 (Z[13], n_220, n_92);
  xnor g188 (Z[14], n_222, n_102);
  xnor g191 (Z[15], n_225, n_98);
  xnor g193 (Z[16], n_189, n_227);
  not g196 (n_66, A[2]);
  not g197 (n_62, A[3]);
  not g198 (n_72, A[4]);
  not g199 (n_68, A[5]);
  not g200 (n_78, A[6]);
  not g201 (n_74, A[7]);
  not g202 (n_84, A[8]);
  not g203 (n_80, A[9]);
  not g204 (n_90, A[10]);
  not g205 (n_86, A[11]);
  not g206 (n_96, A[12]);
  not g207 (n_92, A[13]);
  not g208 (n_102, A[14]);
  not g209 (n_98, A[15]);
  not g211 (n_57, n_37);
  not g212 (n_193, A[1]);
  not g213 (n_227, A[16]);
  not g214 (n_103, n_60);
  not g215 (n_196, n_105);
  not g216 (n_139, n_108);
  not g217 (n_200, n_141);
  not g218 (n_202, n_142);
  not g219 (n_205, n_146);
  not g220 (n_166, n_150);
  not g221 (n_209, n_168);
  not g222 (n_211, n_169);
  not g223 (n_214, n_173);
  not g224 (n_217, n_175);
  not g225 (n_220, n_178);
  not g226 (n_222, n_181);
  not g227 (n_225, n_184);
  not g228 (n_189, n_187);
endmodule

module fx68k_sub_unsigned_1875(A, B, Z);
  input [15:0] A, B;
  output [16:0] Z;
  wire [15:0] A, B;
  wire [16:0] Z;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237;
  not g2 (n_52, B[15]);
  not g3 (n_53, B[14]);
  not g4 (n_54, B[13]);
  not g5 (n_55, B[12]);
  not g6 (n_56, B[11]);
  not g7 (n_57, B[10]);
  not g8 (n_58, B[9]);
  not g9 (n_59, B[8]);
  not g10 (n_60, B[7]);
  not g11 (n_61, B[6]);
  not g12 (n_62, B[5]);
  not g13 (n_63, B[4]);
  not g14 (n_64, B[3]);
  not g15 (n_65, B[2]);
  not g16 (n_66, B[1]);
  not g17 (n_67, B[0]);
  not g18 (Z[16], n_68);
  xor g19 (n_237, A[0], n_67);
  nand g22 (n_72, n_69, B[0]);
  nor g23 (n_71, A[1], n_66);
  nand g24 (n_74, A[1], n_66);
  nor g25 (n_81, A[2], n_65);
  nand g26 (n_76, A[2], n_65);
  nor g27 (n_77, A[3], n_64);
  nand g28 (n_78, A[3], n_64);
  nor g29 (n_87, A[4], n_63);
  nand g30 (n_82, A[4], n_63);
  nor g31 (n_83, A[5], n_62);
  nand g32 (n_84, A[5], n_62);
  nor g33 (n_93, A[6], n_61);
  nand g34 (n_88, A[6], n_61);
  nor g35 (n_89, A[7], n_60);
  nand g36 (n_90, A[7], n_60);
  nor g37 (n_99, A[8], n_59);
  nand g38 (n_94, A[8], n_59);
  nor g39 (n_95, A[9], n_58);
  nand g40 (n_96, A[9], n_58);
  nor g41 (n_105, A[10], n_57);
  nand g42 (n_100, A[10], n_57);
  nor g43 (n_101, A[11], n_56);
  nand g44 (n_102, A[11], n_56);
  nor g45 (n_111, A[12], n_55);
  nand g46 (n_106, A[12], n_55);
  nor g47 (n_107, A[13], n_54);
  nand g48 (n_108, A[13], n_54);
  nor g49 (n_117, A[14], n_53);
  nand g50 (n_112, A[14], n_53);
  nor g51 (n_113, A[15], n_52);
  nand g52 (n_114, A[15], n_52);
  not g53 (n_73, n_71);
  nand g54 (n_75, n_72, n_73);
  nand g55 (n_118, n_74, n_75);
  nor g56 (n_79, n_76, n_77);
  not g57 (n_80, n_78);
  nor g58 (n_122, n_79, n_80);
  nor g59 (n_121, n_81, n_77);
  nor g60 (n_85, n_82, n_83);
  not g61 (n_86, n_84);
  nor g62 (n_124, n_85, n_86);
  nor g63 (n_127, n_87, n_83);
  nor g64 (n_91, n_88, n_89);
  not g65 (n_92, n_90);
  nor g66 (n_131, n_91, n_92);
  nor g67 (n_129, n_93, n_89);
  nor g68 (n_97, n_94, n_95);
  not g69 (n_98, n_96);
  nor g70 (n_134, n_97, n_98);
  nor g71 (n_137, n_99, n_95);
  nor g72 (n_103, n_100, n_101);
  not g73 (n_104, n_102);
  nor g74 (n_141, n_103, n_104);
  nor g75 (n_139, n_105, n_101);
  nor g76 (n_109, n_106, n_107);
  not g77 (n_110, n_108);
  nor g78 (n_144, n_109, n_110);
  nor g79 (n_147, n_111, n_107);
  nor g80 (n_115, n_112, n_113);
  not g81 (n_116, n_114);
  nor g82 (n_151, n_115, n_116);
  nor g83 (n_149, n_117, n_113);
  not g84 (n_119, n_81);
  nand g85 (n_120, n_118, n_119);
  nand g86 (n_206, n_76, n_120);
  nand g87 (n_123, n_121, n_118);
  nand g88 (n_154, n_122, n_123);
  nor g89 (n_125, n_93, n_124);
  not g90 (n_126, n_88);
  nor g91 (n_160, n_125, n_126);
  not g92 (n_128, n_93);
  nand g93 (n_158, n_127, n_128);
  not g94 (n_130, n_129);
  nor g95 (n_132, n_124, n_130);
  not g96 (n_133, n_131);
  nor g97 (n_164, n_132, n_133);
  nand g98 (n_162, n_127, n_129);
  nor g99 (n_135, n_105, n_134);
  not g100 (n_136, n_100);
  nor g101 (n_187, n_135, n_136);
  not g102 (n_138, n_105);
  nand g103 (n_185, n_137, n_138);
  not g104 (n_140, n_139);
  nor g105 (n_142, n_134, n_140);
  not g106 (n_143, n_141);
  nor g107 (n_166, n_142, n_143);
  nand g108 (n_169, n_137, n_139);
  nor g109 (n_145, n_117, n_144);
  not g110 (n_146, n_112);
  nor g111 (n_174, n_145, n_146);
  not g112 (n_148, n_117);
  nand g113 (n_173, n_147, n_148);
  not g114 (n_150, n_149);
  nor g115 (n_152, n_144, n_150);
  not g116 (n_153, n_151);
  nor g117 (n_178, n_152, n_153);
  nand g118 (n_177, n_147, n_149);
  not g119 (n_155, n_87);
  nand g120 (n_156, n_154, n_155);
  nand g121 (n_210, n_82, n_156);
  nand g122 (n_157, n_127, n_154);
  nand g123 (n_212, n_124, n_157);
  not g124 (n_159, n_158);
  nand g125 (n_161, n_154, n_159);
  nand g126 (n_215, n_160, n_161);
  not g127 (n_163, n_162);
  nand g128 (n_165, n_154, n_163);
  nand g129 (n_181, n_164, n_165);
  nor g130 (n_167, n_111, n_166);
  not g131 (n_168, n_106);
  nor g132 (n_192, n_167, n_168);
  nor g133 (n_191, n_111, n_169);
  not g134 (n_170, n_147);
  nor g135 (n_171, n_166, n_170);
  not g136 (n_172, n_144);
  nor g137 (n_195, n_171, n_172);
  nor g138 (n_194, n_169, n_170);
  nor g139 (n_175, n_173, n_166);
  not g140 (n_176, n_174);
  nor g141 (n_198, n_175, n_176);
  nor g142 (n_197, n_169, n_173);
  nor g143 (n_179, n_177, n_166);
  not g144 (n_180, n_178);
  nor g145 (n_201, n_179, n_180);
  nor g146 (n_200, n_169, n_177);
  not g147 (n_182, n_99);
  nand g148 (n_183, n_181, n_182);
  nand g149 (n_219, n_94, n_183);
  nand g150 (n_184, n_137, n_181);
  nand g151 (n_221, n_134, n_184);
  not g152 (n_186, n_185);
  nand g153 (n_188, n_181, n_186);
  nand g154 (n_224, n_187, n_188);
  not g155 (n_189, n_169);
  nand g156 (n_190, n_181, n_189);
  nand g157 (n_227, n_166, n_190);
  nand g158 (n_193, n_191, n_181);
  nand g159 (n_230, n_192, n_193);
  nand g160 (n_196, n_194, n_181);
  nand g161 (n_232, n_195, n_196);
  nand g162 (n_199, n_197, n_181);
  nand g163 (n_235, n_198, n_199);
  nand g164 (n_202, n_200, n_181);
  nand g165 (n_68, n_201, n_202);
  nand g166 (n_203, n_73, n_74);
  xnor g167 (Z[1], n_72, n_203);
  nand g168 (n_204, n_119, n_76);
  xnor g169 (Z[2], n_118, n_204);
  not g170 (n_205, n_77);
  nand g171 (n_207, n_205, n_78);
  xnor g172 (Z[3], n_206, n_207);
  nand g173 (n_208, n_155, n_82);
  xnor g174 (Z[4], n_154, n_208);
  not g175 (n_209, n_83);
  nand g176 (n_211, n_209, n_84);
  xnor g177 (Z[5], n_210, n_211);
  nand g178 (n_213, n_128, n_88);
  xnor g179 (Z[6], n_212, n_213);
  not g180 (n_214, n_89);
  nand g181 (n_216, n_214, n_90);
  xnor g182 (Z[7], n_215, n_216);
  nand g183 (n_217, n_182, n_94);
  xnor g184 (Z[8], n_181, n_217);
  not g185 (n_218, n_95);
  nand g186 (n_220, n_218, n_96);
  xnor g187 (Z[9], n_219, n_220);
  nand g188 (n_222, n_138, n_100);
  xnor g189 (Z[10], n_221, n_222);
  not g190 (n_223, n_101);
  nand g191 (n_225, n_223, n_102);
  xnor g192 (Z[11], n_224, n_225);
  not g193 (n_226, n_111);
  nand g194 (n_228, n_226, n_106);
  xnor g195 (Z[12], n_227, n_228);
  not g196 (n_229, n_107);
  nand g197 (n_231, n_229, n_108);
  xnor g198 (Z[13], n_230, n_231);
  nand g199 (n_233, n_148, n_112);
  xnor g200 (Z[14], n_232, n_233);
  not g201 (n_234, n_113);
  nand g202 (n_236, n_234, n_114);
  xnor g203 (Z[15], n_235, n_236);
  not g205 (n_69, A[0]);
  not g206 (Z[0], n_237);
endmodule

module fx68k_sub_signed_1877(A, B, Z);
  input [16:0] A;
  input [1:0] B;
  output [16:0] Z;
  wire [16:0] A;
  wire [1:0] B;
  wire [16:0] Z;
  wire n_39, n_40, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_73, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  not g2 (n_39, B[0]);
  not g3 (n_40, B[1]);
  not g18 (n_55, A[16]);
  xor g20 (n_232, A[0], n_39);
  nand g23 (n_76, n_73, B[0]);
  nor g24 (n_75, A[1], n_40);
  nand g25 (n_78, A[1], n_40);
  nor g26 (n_85, A[2], n_40);
  nand g27 (n_80, A[2], n_40);
  nor g28 (n_81, A[3], n_40);
  nand g29 (n_82, A[3], n_40);
  nor g30 (n_91, A[4], n_40);
  nand g31 (n_86, A[4], n_40);
  nor g32 (n_87, A[5], n_40);
  nand g33 (n_88, A[5], n_40);
  nor g34 (n_60, A[6], n_40);
  nand g35 (n_92, A[6], n_40);
  nor g36 (n_56, A[7], n_40);
  nand g37 (n_57, A[7], n_40);
  nor g38 (n_66, A[8], n_40);
  nand g39 (n_61, A[8], n_40);
  nor g40 (n_62, A[9], n_40);
  nand g41 (n_63, A[9], n_40);
  nor g42 (n_94, A[10], n_40);
  nand g43 (n_67, A[10], n_40);
  nor g44 (n_68, A[11], n_40);
  nand g45 (n_69, A[11], n_40);
  nor g46 (n_100, A[12], n_40);
  nand g47 (n_95, A[12], n_40);
  nor g48 (n_96, A[13], n_40);
  nand g49 (n_97, A[13], n_40);
  nor g50 (n_106, A[14], n_40);
  nand g51 (n_101, A[14], n_40);
  nor g52 (n_102, A[15], n_40);
  nand g53 (n_103, A[15], n_40);
  nor g54 (n_192, n_55, B[1]);
  nand g55 (n_195, n_55, B[1]);
  not g56 (n_77, n_75);
  nand g57 (n_79, n_76, n_77);
  nand g58 (n_107, n_78, n_79);
  nor g59 (n_83, n_80, n_81);
  not g60 (n_84, n_82);
  nor g61 (n_111, n_83, n_84);
  nor g62 (n_110, n_85, n_81);
  nor g63 (n_89, n_86, n_87);
  not g64 (n_90, n_88);
  nor g65 (n_113, n_89, n_90);
  nor g66 (n_116, n_91, n_87);
  nor g67 (n_58, n_92, n_56);
  not g68 (n_59, n_57);
  nor g69 (n_120, n_58, n_59);
  nor g70 (n_118, n_60, n_56);
  nor g71 (n_64, n_61, n_62);
  not g72 (n_65, n_63);
  nor g73 (n_123, n_64, n_65);
  nor g74 (n_126, n_66, n_62);
  nor g75 (n_70, n_67, n_68);
  not g76 (n_93, n_69);
  nor g77 (n_130, n_70, n_93);
  nor g78 (n_128, n_94, n_68);
  nor g79 (n_98, n_95, n_96);
  not g80 (n_99, n_97);
  nor g81 (n_133, n_98, n_99);
  nor g82 (n_136, n_100, n_96);
  nor g83 (n_104, n_101, n_102);
  not g84 (n_105, n_103);
  nor g85 (n_140, n_104, n_105);
  nor g86 (n_138, n_106, n_102);
  not g87 (n_108, n_85);
  nand g88 (n_109, n_107, n_108);
  nand g89 (n_200, n_80, n_109);
  nand g90 (n_112, n_110, n_107);
  nand g91 (n_143, n_111, n_112);
  nor g92 (n_114, n_60, n_113);
  not g93 (n_115, n_92);
  nor g94 (n_149, n_114, n_115);
  not g95 (n_117, n_60);
  nand g96 (n_147, n_116, n_117);
  not g97 (n_119, n_118);
  nor g98 (n_121, n_113, n_119);
  not g99 (n_122, n_120);
  nor g100 (n_153, n_121, n_122);
  nand g101 (n_151, n_116, n_118);
  nor g102 (n_124, n_94, n_123);
  not g103 (n_125, n_67);
  nor g104 (n_176, n_124, n_125);
  not g105 (n_127, n_94);
  nand g106 (n_174, n_126, n_127);
  not g107 (n_129, n_128);
  nor g108 (n_131, n_123, n_129);
  not g109 (n_132, n_130);
  nor g110 (n_155, n_131, n_132);
  nand g111 (n_158, n_126, n_128);
  nor g112 (n_134, n_106, n_133);
  not g113 (n_135, n_101);
  nor g114 (n_163, n_134, n_135);
  not g115 (n_137, n_106);
  nand g116 (n_162, n_136, n_137);
  not g117 (n_139, n_138);
  nor g118 (n_141, n_133, n_139);
  not g119 (n_142, n_140);
  nor g120 (n_167, n_141, n_142);
  nand g121 (n_166, n_136, n_138);
  not g122 (n_144, n_91);
  nand g123 (n_145, n_143, n_144);
  nand g124 (n_204, n_86, n_145);
  nand g125 (n_146, n_116, n_143);
  nand g126 (n_206, n_113, n_146);
  not g127 (n_148, n_147);
  nand g128 (n_150, n_143, n_148);
  nand g129 (n_209, n_149, n_150);
  not g130 (n_152, n_151);
  nand g131 (n_154, n_143, n_152);
  nand g132 (n_170, n_153, n_154);
  nor g133 (n_156, n_100, n_155);
  not g134 (n_157, n_95);
  nor g135 (n_181, n_156, n_157);
  nor g136 (n_180, n_100, n_158);
  not g137 (n_159, n_136);
  nor g138 (n_160, n_155, n_159);
  not g139 (n_161, n_133);
  nor g140 (n_184, n_160, n_161);
  nor g141 (n_183, n_158, n_159);
  nor g142 (n_164, n_162, n_155);
  not g143 (n_165, n_163);
  nor g144 (n_187, n_164, n_165);
  nor g145 (n_186, n_158, n_162);
  nor g146 (n_168, n_166, n_155);
  not g147 (n_169, n_167);
  nor g148 (n_190, n_168, n_169);
  nor g149 (n_189, n_158, n_166);
  not g150 (n_171, n_66);
  nand g151 (n_172, n_170, n_171);
  nand g152 (n_213, n_61, n_172);
  nand g153 (n_173, n_126, n_170);
  nand g154 (n_215, n_123, n_173);
  not g155 (n_175, n_174);
  nand g156 (n_177, n_170, n_175);
  nand g157 (n_218, n_176, n_177);
  not g158 (n_178, n_158);
  nand g159 (n_179, n_170, n_178);
  nand g160 (n_221, n_155, n_179);
  nand g161 (n_182, n_180, n_170);
  nand g162 (n_224, n_181, n_182);
  nand g163 (n_185, n_183, n_170);
  nand g164 (n_226, n_184, n_185);
  nand g165 (n_188, n_186, n_170);
  nand g166 (n_229, n_187, n_188);
  nand g167 (n_191, n_189, n_170);
  nand g168 (n_193, n_190, n_191);
  not g169 (n_194, n_192);
  nand g172 (n_197, n_77, n_78);
  xnor g173 (Z[1], n_76, n_197);
  nand g174 (n_198, n_108, n_80);
  xnor g175 (Z[2], n_107, n_198);
  not g176 (n_199, n_81);
  nand g177 (n_201, n_199, n_82);
  xnor g178 (Z[3], n_200, n_201);
  nand g179 (n_202, n_144, n_86);
  xnor g180 (Z[4], n_143, n_202);
  not g181 (n_203, n_87);
  nand g182 (n_205, n_203, n_88);
  xnor g183 (Z[5], n_204, n_205);
  nand g184 (n_207, n_117, n_92);
  xnor g185 (Z[6], n_206, n_207);
  not g186 (n_208, n_56);
  nand g187 (n_210, n_208, n_57);
  xnor g188 (Z[7], n_209, n_210);
  nand g189 (n_211, n_171, n_61);
  xnor g190 (Z[8], n_170, n_211);
  not g191 (n_212, n_62);
  nand g192 (n_214, n_212, n_63);
  xnor g193 (Z[9], n_213, n_214);
  nand g194 (n_216, n_127, n_67);
  xnor g195 (Z[10], n_215, n_216);
  not g196 (n_217, n_68);
  nand g197 (n_219, n_217, n_69);
  xnor g198 (Z[11], n_218, n_219);
  not g199 (n_220, n_100);
  nand g200 (n_222, n_220, n_95);
  xnor g201 (Z[12], n_221, n_222);
  not g202 (n_223, n_96);
  nand g203 (n_225, n_223, n_97);
  xnor g204 (Z[13], n_224, n_225);
  nand g205 (n_227, n_137, n_101);
  xnor g206 (Z[14], n_226, n_227);
  not g207 (n_228, n_102);
  nand g208 (n_230, n_228, n_103);
  xnor g209 (Z[15], n_229, n_230);
  nand g210 (n_231, n_194, n_195);
  xnor g211 (Z[16], n_193, n_231);
  not g213 (n_73, A[0]);
  not g214 (Z[0], n_232);
endmodule

module fx68k_bmux_1882(ctl, in_0, in_1, z);
  input ctl;
  input [15:0] in_0, in_1;
  output [15:0] z;
  wire ctl;
  wire [15:0] in_0, in_1;
  wire [15:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[15]), .data1 (in_1[15]), .z
       (z[15]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[14]), .data1 (in_1[14]), .z
       (z[14]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[13]), .data1 (in_1[13]), .z
       (z[13]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[12]), .data1 (in_1[12]), .z
       (z[12]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[11]), .data1 (in_1[11]), .z
       (z[11]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[10]), .data1 (in_1[10]), .z
       (z[10]));
  CDN_bmux2 g7(.sel0 (ctl), .data0 (in_0[9]), .data1 (in_1[9]), .z
       (z[9]));
  CDN_bmux2 g8(.sel0 (ctl), .data0 (in_0[8]), .data1 (in_1[8]), .z
       (z[8]));
  CDN_bmux2 g9(.sel0 (ctl), .data0 (in_0[7]), .data1 (in_1[7]), .z
       (z[7]));
  CDN_bmux2 g10(.sel0 (ctl), .data0 (in_0[6]), .data1 (in_1[6]), .z
       (z[6]));
  CDN_bmux2 g11(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g12(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g13(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g14(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g15(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g16(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_bmux_1883(ctl, in_0, in_1, in_2, in_3, z);
  input [1:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3;
  output [15:0] z;
  wire [1:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3;
  wire [15:0] z;
  CDN_bmux4 g1(.sel0 (ctl[0]), .data0 (in_0[15]), .data1 (in_1[15]),
       .sel1 (ctl[1]), .data2 (in_2[15]), .data3 (in_3[15]), .z
       (z[15]));
  CDN_bmux4 g2(.sel0 (ctl[0]), .data0 (in_0[14]), .data1 (in_1[14]),
       .sel1 (ctl[1]), .data2 (in_2[14]), .data3 (in_3[14]), .z
       (z[14]));
  CDN_bmux4 g3(.sel0 (ctl[0]), .data0 (in_0[13]), .data1 (in_1[13]),
       .sel1 (ctl[1]), .data2 (in_2[13]), .data3 (in_3[13]), .z
       (z[13]));
  CDN_bmux4 g4(.sel0 (ctl[0]), .data0 (in_0[12]), .data1 (in_1[12]),
       .sel1 (ctl[1]), .data2 (in_2[12]), .data3 (in_3[12]), .z
       (z[12]));
  CDN_bmux4 g5(.sel0 (ctl[0]), .data0 (in_0[11]), .data1 (in_1[11]),
       .sel1 (ctl[1]), .data2 (in_2[11]), .data3 (in_3[11]), .z
       (z[11]));
  CDN_bmux4 g6(.sel0 (ctl[0]), .data0 (in_0[10]), .data1 (in_1[10]),
       .sel1 (ctl[1]), .data2 (in_2[10]), .data3 (in_3[10]), .z
       (z[10]));
  CDN_bmux4 g7(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .z (z[9]));
  CDN_bmux4 g8(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .z (z[8]));
  CDN_bmux4 g9(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .z (z[7]));
  CDN_bmux4 g10(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .z (z[6]));
  CDN_bmux4 g11(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .z (z[5]));
  CDN_bmux4 g12(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .z (z[4]));
  CDN_bmux4 g13(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .z (z[3]));
  CDN_bmux4 g14(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .z (z[2]));
  CDN_bmux4 g15(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .z (z[1]));
  CDN_bmux4 g16(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_case_box_1144(in_0, out_0);
  input [4:0] in_0;
  output [9:0] out_0;
  wire [4:0] in_0;
  wire [9:0] out_0;
  wire n_6, n_7, n_8, n_13, n_20, n_31, n_34, n_48;
  wire n_73, n_74, n_75, n_76, n_106, n_107;
  nand g1 (n_6, in_0[4], n_106, in_0[2], n_107);
  not g2 (n_7, in_0[0]);
  nor g3 (out_0[9], n_6, n_7);
  nand g4 (n_13, n_8, in_0[3], in_0[2], n_107);
  nor g6 (out_0[8], n_13, n_7);
  nand g7 (n_20, n_8, in_0[3], in_0[2], in_0[1]);
  nor g9 (out_0[7], n_20, in_0[0]);
  nor g12 (out_0[6], n_20, n_7);
  nand g13 (n_34, in_0[4], n_106, n_31, n_107);
  nor g15 (out_0[5], n_34, in_0[0]);
  nor g18 (out_0[4], n_34, n_7);
  nand g19 (n_48, in_0[4], n_106, n_31, in_0[1]);
  nor g21 (out_0[3], n_48, in_0[0]);
  nor g24 (out_0[2], n_48, n_7);
  nor g27 (out_0[1], n_6, in_0[0]);
  nor g28 (n_74, out_0[9], out_0[8], out_0[7], out_0[6]);
  nor g29 (n_75, out_0[5], out_0[4], out_0[3], out_0[2]);
  not g30 (n_73, out_0[1]);
  nand g31 (n_76, n_73, n_74, n_75);
  not g32 (out_0[0], n_76);
  not g33 (n_106, in_0[3]);
  not g34 (n_107, in_0[1]);
  not g35 (n_8, in_0[4]);
  not g36 (n_31, in_0[2]);
endmodule

module fx68k_mux_1884(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, z);
  input [9:0] ctl;
  input [1:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9;
  output [1:0] z;
  wire [9:0] ctl;
  wire [1:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9;
  wire [1:0] z;
  CDN_mux10 g1(.sel0 (ctl[9]), .data0 (in_0[1]), .sel1 (ctl[8]), .data1
       (in_1[1]), .sel2 (ctl[7]), .data2 (in_2[1]), .sel3 (ctl[6]),
       .data3 (in_3[1]), .sel4 (ctl[5]), .data4 (in_4[1]), .sel5
       (ctl[4]), .data5 (in_5[1]), .sel6 (ctl[3]), .data6 (in_6[1]),
       .sel7 (ctl[2]), .data7 (in_7[1]), .sel8 (ctl[1]), .data8
       (in_8[1]), .sel9 (ctl[0]), .data9 (in_9[1]), .z (z[1]));
  CDN_mux10 g3(.sel0 (ctl[9]), .data0 (in_0[0]), .sel1 (ctl[8]), .data1
       (in_1[0]), .sel2 (ctl[7]), .data2 (in_2[0]), .sel3 (ctl[6]),
       .data3 (in_3[0]), .sel4 (ctl[5]), .data4 (in_4[0]), .sel5
       (ctl[4]), .data5 (in_5[0]), .sel6 (ctl[3]), .data6 (in_6[0]),
       .sel7 (ctl[2]), .data7 (in_7[0]), .sel8 (ctl[1]), .data8
       (in_8[0]), .sel9 (ctl[0]), .data9 (in_9[0]), .z (z[0]));
endmodule

module fx68k_bmux_1894(ctl, in_0, in_1, z);
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[16]), .data1 (in_1[16]), .z
       (z[16]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[15]), .data1 (in_1[15]), .z
       (z[15]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[14]), .data1 (in_1[14]), .z
       (z[14]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[13]), .data1 (in_1[13]), .z
       (z[13]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[12]), .data1 (in_1[12]), .z
       (z[12]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[11]), .data1 (in_1[11]), .z
       (z[11]));
  CDN_bmux2 g7(.sel0 (ctl), .data0 (in_0[10]), .data1 (in_1[10]), .z
       (z[10]));
  CDN_bmux2 g8(.sel0 (ctl), .data0 (in_0[9]), .data1 (in_1[9]), .z
       (z[9]));
  CDN_bmux2 g9(.sel0 (ctl), .data0 (in_0[8]), .data1 (in_1[8]), .z
       (z[8]));
  CDN_bmux2 g10(.sel0 (ctl), .data0 (in_0[7]), .data1 (in_1[7]), .z
       (z[7]));
  CDN_bmux2 g11(.sel0 (ctl), .data0 (in_0[6]), .data1 (in_1[6]), .z
       (z[6]));
  CDN_bmux2 g12(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g13(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g14(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g15(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g16(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g17(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k_mux_1906(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output [15:0] z;
  wire [6:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire [15:0] z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0[15]), .sel1 (ctl[5]), .data1
       (in_1[15]), .sel2 (ctl[4]), .data2 (in_2[15]), .sel3 (ctl[3]),
       .data3 (in_3[15]), .sel4 (ctl[2]), .data4 (in_4[15]), .sel5
       (ctl[1]), .data5 (in_5[15]), .sel6 (ctl[0]), .data6 (in_6[15]),
       .z (z[15]));
  CDN_mux7 g17(.sel0 (ctl[6]), .data0 (in_0[14]), .sel1 (ctl[5]),
       .data1 (in_1[14]), .sel2 (ctl[4]), .data2 (in_2[14]), .sel3
       (ctl[3]), .data3 (in_3[14]), .sel4 (ctl[2]), .data4 (in_4[14]),
       .sel5 (ctl[1]), .data5 (in_5[14]), .sel6 (ctl[0]), .data6
       (in_6[14]), .z (z[14]));
  CDN_mux7 g18(.sel0 (ctl[6]), .data0 (in_0[13]), .sel1 (ctl[5]),
       .data1 (in_1[13]), .sel2 (ctl[4]), .data2 (in_2[13]), .sel3
       (ctl[3]), .data3 (in_3[13]), .sel4 (ctl[2]), .data4 (in_4[13]),
       .sel5 (ctl[1]), .data5 (in_5[13]), .sel6 (ctl[0]), .data6
       (in_6[13]), .z (z[13]));
  CDN_mux7 g19(.sel0 (ctl[6]), .data0 (in_0[12]), .sel1 (ctl[5]),
       .data1 (in_1[12]), .sel2 (ctl[4]), .data2 (in_2[12]), .sel3
       (ctl[3]), .data3 (in_3[12]), .sel4 (ctl[2]), .data4 (in_4[12]),
       .sel5 (ctl[1]), .data5 (in_5[12]), .sel6 (ctl[0]), .data6
       (in_6[12]), .z (z[12]));
  CDN_mux7 g20(.sel0 (ctl[6]), .data0 (in_0[11]), .sel1 (ctl[5]),
       .data1 (in_1[11]), .sel2 (ctl[4]), .data2 (in_2[11]), .sel3
       (ctl[3]), .data3 (in_3[11]), .sel4 (ctl[2]), .data4 (in_4[11]),
       .sel5 (ctl[1]), .data5 (in_5[11]), .sel6 (ctl[0]), .data6
       (in_6[11]), .z (z[11]));
  CDN_mux7 g21(.sel0 (ctl[6]), .data0 (in_0[10]), .sel1 (ctl[5]),
       .data1 (in_1[10]), .sel2 (ctl[4]), .data2 (in_2[10]), .sel3
       (ctl[3]), .data3 (in_3[10]), .sel4 (ctl[2]), .data4 (in_4[10]),
       .sel5 (ctl[1]), .data5 (in_5[10]), .sel6 (ctl[0]), .data6
       (in_6[10]), .z (z[10]));
  CDN_mux7 g22(.sel0 (ctl[6]), .data0 (in_0[9]), .sel1 (ctl[5]), .data1
       (in_1[9]), .sel2 (ctl[4]), .data2 (in_2[9]), .sel3 (ctl[3]),
       .data3 (in_3[9]), .sel4 (ctl[2]), .data4 (in_4[9]), .sel5
       (ctl[1]), .data5 (in_5[9]), .sel6 (ctl[0]), .data6 (in_6[9]), .z
       (z[9]));
  CDN_mux7 g23(.sel0 (ctl[6]), .data0 (in_0[8]), .sel1 (ctl[5]), .data1
       (in_1[8]), .sel2 (ctl[4]), .data2 (in_2[8]), .sel3 (ctl[3]),
       .data3 (in_3[8]), .sel4 (ctl[2]), .data4 (in_4[8]), .sel5
       (ctl[1]), .data5 (in_5[8]), .sel6 (ctl[0]), .data6 (in_6[8]), .z
       (z[8]));
  CDN_mux7 g24(.sel0 (ctl[6]), .data0 (in_0[7]), .sel1 (ctl[5]), .data1
       (in_1[7]), .sel2 (ctl[4]), .data2 (in_2[7]), .sel3 (ctl[3]),
       .data3 (in_3[7]), .sel4 (ctl[2]), .data4 (in_4[7]), .sel5
       (ctl[1]), .data5 (in_5[7]), .sel6 (ctl[0]), .data6 (in_6[7]), .z
       (z[7]));
  CDN_mux7 g25(.sel0 (ctl[6]), .data0 (in_0[6]), .sel1 (ctl[5]), .data1
       (in_1[6]), .sel2 (ctl[4]), .data2 (in_2[6]), .sel3 (ctl[3]),
       .data3 (in_3[6]), .sel4 (ctl[2]), .data4 (in_4[6]), .sel5
       (ctl[1]), .data5 (in_5[6]), .sel6 (ctl[0]), .data6 (in_6[6]), .z
       (z[6]));
  CDN_mux7 g26(.sel0 (ctl[6]), .data0 (in_0[5]), .sel1 (ctl[5]), .data1
       (in_1[5]), .sel2 (ctl[4]), .data2 (in_2[5]), .sel3 (ctl[3]),
       .data3 (in_3[5]), .sel4 (ctl[2]), .data4 (in_4[5]), .sel5
       (ctl[1]), .data5 (in_5[5]), .sel6 (ctl[0]), .data6 (in_6[5]), .z
       (z[5]));
  CDN_mux7 g27(.sel0 (ctl[6]), .data0 (in_0[4]), .sel1 (ctl[5]), .data1
       (in_1[4]), .sel2 (ctl[4]), .data2 (in_2[4]), .sel3 (ctl[3]),
       .data3 (in_3[4]), .sel4 (ctl[2]), .data4 (in_4[4]), .sel5
       (ctl[1]), .data5 (in_5[4]), .sel6 (ctl[0]), .data6 (in_6[4]), .z
       (z[4]));
  CDN_mux7 g28(.sel0 (ctl[6]), .data0 (in_0[3]), .sel1 (ctl[5]), .data1
       (in_1[3]), .sel2 (ctl[4]), .data2 (in_2[3]), .sel3 (ctl[3]),
       .data3 (in_3[3]), .sel4 (ctl[2]), .data4 (in_4[3]), .sel5
       (ctl[1]), .data5 (in_5[3]), .sel6 (ctl[0]), .data6 (in_6[3]), .z
       (z[3]));
  CDN_mux7 g29(.sel0 (ctl[6]), .data0 (in_0[2]), .sel1 (ctl[5]), .data1
       (in_1[2]), .sel2 (ctl[4]), .data2 (in_2[2]), .sel3 (ctl[3]),
       .data3 (in_3[2]), .sel4 (ctl[2]), .data4 (in_4[2]), .sel5
       (ctl[1]), .data5 (in_5[2]), .sel6 (ctl[0]), .data6 (in_6[2]), .z
       (z[2]));
  CDN_mux7 g30(.sel0 (ctl[6]), .data0 (in_0[1]), .sel1 (ctl[5]), .data1
       (in_1[1]), .sel2 (ctl[4]), .data2 (in_2[1]), .sel3 (ctl[3]),
       .data3 (in_3[1]), .sel4 (ctl[2]), .data4 (in_4[1]), .sel5
       (ctl[1]), .data5 (in_5[1]), .sel6 (ctl[0]), .data6 (in_6[1]), .z
       (z[1]));
  CDN_mux7 g31(.sel0 (ctl[6]), .data0 (in_0[0]), .sel1 (ctl[5]), .data1
       (in_1[0]), .sel2 (ctl[4]), .data2 (in_2[0]), .sel3 (ctl[3]),
       .data3 (in_3[0]), .sel4 (ctl[2]), .data4 (in_4[0]), .sel5
       (ctl[1]), .data5 (in_5[0]), .sel6 (ctl[0]), .data6 (in_6[0]), .z
       (z[0]));
endmodule

module fx68k_mux_1926(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, z);
  input [11:0] ctl;
  input [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  output [3:0] z;
  wire [11:0] ctl;
  wire [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11;
  wire [3:0] z;
  CDN_mux12 g1(.sel0 (ctl[11]), .data0 (in_0[3]), .sel1 (ctl[10]),
       .data1 (in_1[3]), .sel2 (ctl[9]), .data2 (in_2[3]), .sel3
       (ctl[8]), .data3 (in_3[3]), .sel4 (ctl[7]), .data4 (in_4[3]),
       .sel5 (ctl[6]), .data5 (in_5[3]), .sel6 (ctl[5]), .data6
       (in_6[3]), .sel7 (ctl[4]), .data7 (in_7[3]), .sel8 (ctl[3]),
       .data8 (in_8[3]), .sel9 (ctl[2]), .data9 (in_9[3]), .sel10
       (ctl[1]), .data10 (in_10[3]), .sel11 (ctl[0]), .data11
       (in_11[3]), .z (z[3]));
  CDN_mux12 g5(.sel0 (ctl[11]), .data0 (in_0[2]), .sel1 (ctl[10]),
       .data1 (in_1[2]), .sel2 (ctl[9]), .data2 (in_2[2]), .sel3
       (ctl[8]), .data3 (in_3[2]), .sel4 (ctl[7]), .data4 (in_4[2]),
       .sel5 (ctl[6]), .data5 (in_5[2]), .sel6 (ctl[5]), .data6
       (in_6[2]), .sel7 (ctl[4]), .data7 (in_7[2]), .sel8 (ctl[3]),
       .data8 (in_8[2]), .sel9 (ctl[2]), .data9 (in_9[2]), .sel10
       (ctl[1]), .data10 (in_10[2]), .sel11 (ctl[0]), .data11
       (in_11[2]), .z (z[2]));
  CDN_mux12 g6(.sel0 (ctl[11]), .data0 (in_0[1]), .sel1 (ctl[10]),
       .data1 (in_1[1]), .sel2 (ctl[9]), .data2 (in_2[1]), .sel3
       (ctl[8]), .data3 (in_3[1]), .sel4 (ctl[7]), .data4 (in_4[1]),
       .sel5 (ctl[6]), .data5 (in_5[1]), .sel6 (ctl[5]), .data6
       (in_6[1]), .sel7 (ctl[4]), .data7 (in_7[1]), .sel8 (ctl[3]),
       .data8 (in_8[1]), .sel9 (ctl[2]), .data9 (in_9[1]), .sel10
       (ctl[1]), .data10 (in_10[1]), .sel11 (ctl[0]), .data11
       (in_11[1]), .z (z[1]));
  CDN_mux12 g7(.sel0 (ctl[11]), .data0 (in_0[0]), .sel1 (ctl[10]),
       .data1 (in_1[0]), .sel2 (ctl[9]), .data2 (in_2[0]), .sel3
       (ctl[8]), .data3 (in_3[0]), .sel4 (ctl[7]), .data4 (in_4[0]),
       .sel5 (ctl[6]), .data5 (in_5[0]), .sel6 (ctl[5]), .data6
       (in_6[0]), .sel7 (ctl[4]), .data7 (in_7[0]), .sel8 (ctl[3]),
       .data8 (in_8[0]), .sel9 (ctl[2]), .data9 (in_9[0]), .sel10
       (ctl[1]), .data10 (in_10[0]), .sel11 (ctl[0]), .data11
       (in_11[0]), .z (z[0]));
endmodule

module fx68k_fx68kAlu(clk, pwrUp, enT1, enT3, enT4, ird, aluColumn,
     aluDataCtrl, aluAddrCtrl, alueClkEn, ftu2Ccr, init, finish,
     aluIsByte, ftu, alub, iDataBus, iAddrBus, ze, alue, ccr, aluOut);
  input clk, pwrUp, enT1, enT3, enT4, aluAddrCtrl, alueClkEn, ftu2Ccr,
       init, finish, aluIsByte;
  input [15:0] ird, ftu, alub, iDataBus, iAddrBus;
  input [2:0] aluColumn;
  input [1:0] aluDataCtrl;
  output ze;
  output [15:0] alue, aluOut;
  output [7:0] ccr;
  wire clk, pwrUp, enT1, enT3, enT4, aluAddrCtrl, alueClkEn, ftu2Ccr,
       init, finish, aluIsByte;
  wire [15:0] ird, ftu, alub, iDataBus, iAddrBus;
  wire [2:0] aluColumn;
  wire [1:0] aluDataCtrl;
  wire ze;
  wire [15:0] alue, aluOut;
  wire [7:0] ccr;
  wire [15:0] cRow;
  wire [15:0] row;
  wire [4:0] aluOp;
  wire [4:0] cMask;
  wire [15:0] aOperand;
  wire [1:0] cmbsop_isShift;
  wire [31:0] shftResult;
  wire [7:0] bcdResult;
  wire [4:0] ccrCore;
  wire [15:0] inpb;
  wire [15:0] result;
  wire [4:0] ccrTemp;
  wire [4:0] ccrMask;
  wire [4:0] ccrMasked;
  wire [16:0] rtemp;
  wire [4:0] oper;
  wire [15:0] mySubber_228_3;
  wire [7:0] bcdLatch;
  wire UNCONNECTED437, UNCONNECTED438, UNCONNECTED439, UNCONNECTED440,
       UNCONNECTED441, _X_, bAdd, bcdC;
  wire bcdCarry, bcdOverf, bcdV, cIsArX, cNoCcrEn, cin, coreH, dm;
  wire isArX, isByte, isCorf, isLong, n_6, n_7, n_8, n_9;
  wire n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17;
  wire n_19, n_20, n_21, n_23, n_24, n_25, n_26, n_27;
  wire n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_36;
  wire n_37, n_38, n_39, n_40, n_42, n_43, n_82, n_98;
  wire n_151, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_165, n_167, n_169, n_170;
  wire n_171, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_226, n_227, n_228, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_404, n_405, n_406, n_407, n_408, n_411, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_464, n_465, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_498, n_499, n_500, n_501, n_502, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_531, n_707, n_708, n_709, n_712;
  wire n_714, n_717, n_718, n_723, n_724, n_730, n_733, n_735;
  wire n_755, n_756, n_757, n_761, n_764, n_766, n_767, n_775;
  wire n_777, n_779, n_780, n_781, n_782, n_783, n_784, n_785;
  wire n_786, n_787, n_788, n_796, n_799, n_800, n_802, n_803;
  wire n_804, n_805, n_806, n_807, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820;
  wire n_822, n_823, n_824, n_825, n_826, noCcrEn, rIrd8, rm;
  wire shftCin, shftMsb, sm, subCout, subHcarry, subOv, tsm;
  assign ccr[5] = 1'b0;
  assign ccr[6] = 1'b0;
  assign ccr[7] = 1'b0;
  fx68k_rowDecoder rowDecoder(.ird (ird), .row (cRow), .noCcrEn
       (cNoCcrEn), .isArX (cIsArX));
  fx68k_aluGetOp aluGetOp(.row (row), .col (aluColumn), .isCorf
       (isCorf), .aluOp (aluOp));
  fx68k_ccrTable ccrTable(.col (aluColumn), .row (row), .finish
       (finish), .ccrMask (cMask));
  fx68k_aluShifter shifter(.data ({alue, aOperand}), .isByte (isByte),
       .isLong (isLong), .swapWords (n_404), .dir (cmbsop_isShift[0]),
       .cin (shftCin), .result (shftResult));
  fx68k_aluCorf aluCorf(.binResult (aluOut[7:0]), .bAdd (n_405), .cin
       (ccr[4]), .hCarry (coreH), .bcdResult (bcdResult), .dC (bcdC),
       .ov (bcdV));
  fx68k_and_op g21(.A (aOperand), .B (inpb), .Z ({n_350, n_347, n_344,
       n_341, n_338, n_335, n_332, n_329, n_326, n_323, n_320, n_317,
       n_314, n_311, n_308, n_305}));
  fx68k_or_op_1132 g22(.A (aOperand), .B (inpb), .Z ({n_351, n_348,
       n_345, n_342, n_339, n_336, n_333, n_330, n_327, n_324, n_321,
       n_318, n_315, n_312, n_309, n_306}));
  fx68k_xor_op g23(.A (aOperand), .B (inpb), .Z ({n_352, n_349, n_346,
       n_343, n_340, n_337, n_334, n_331, n_328, n_325, n_322, n_319,
       n_316, n_313, n_310, n_307}));
  fx68k_or_op_1133 g24(.A (result[7:0]), .Z (n_416));
  fx68k_or_op_1134 g26(.A (result), .Z (n_417));
  fx68k_and_op_1135 g32(.A (ccrTemp), .B (ccrMask), .Z ({n_431, n_430,
       n_429, n_428, n_427}));
  fx68k_not_op g33(.A (ccrMask), .Z ({n_426, n_425, n_424, n_423,
       n_422}));
  fx68k_and_op_1136 g34(.A (ccr[4:0]), .B ({n_426, n_425, n_424, n_423,
       n_422}), .Z ({n_436, n_435, n_434, n_433, n_432}));
  fx68k_or_op_1137 g35(.A ({n_431, n_430, n_429, n_428, n_427}), .B
       ({n_436, n_435, n_434, n_433, n_432}), .Z ({ccrMasked[4:3],
       n_171, ccrMasked[1:0]}));
  fx68k_or_op_1138 g38(.A (aluColumn), .Z (n_98));
  fx68k_add_unsigned_1865 \mySubber_228_3:add_278_39 (.A ({1'b0,
       inpb[7:0]}), .B ({1'b0, aOperand[7:0]}), .Z ({n_486, n_485,
       n_484, n_483, n_482, n_481, n_480, n_479, n_478, n_477}));
  fx68k_add_unsigned_1867 \mySubber_228_3:add_278_60 (.A ({n_486,
       n_485, n_484, n_483, n_482, n_481, n_480, n_479, n_478, n_477}),
       .B (cin), .Z ({n_256, n_254, n_252, n_250, n_248, n_246, n_244,
       n_242, n_240, n_238, n_236}));
  fx68k_sub_unsigned_1869 \mySubber_228_3:sub_279_29 (.A ({1'b0,
       inpb[7:0]}), .B ({1'b0, aOperand[7:0]}), .Z ({n_496, n_495,
       n_494, n_493, n_492, n_491, n_490, n_489, n_488, n_487}));
  fx68k_sub_signed \mySubber_228_3:sub_279_50 (.A ({n_496, n_495,
       n_494, n_493, n_492, n_491, n_490, n_489, n_488, n_487}), .B
       ({1'b0, cin}), .Z ({n_263, n_262, n_261, n_260, n_259, n_258,
       n_257, n_255, n_253, n_251, n_249, n_247, n_245, n_243, n_241,
       n_239, n_237}));
  fx68k_add_unsigned_1871 \mySubber_228_3:add_284_35 (.A (inpb), .B
       (aOperand), .Z ({n_514, n_513, n_512, n_511, n_510, n_509,
       n_508, n_507, n_506, n_505, n_504, n_503, n_502, n_501, n_500,
       n_499, n_498}));
  fx68k_add_unsigned_1873 \mySubber_228_3:add_284_51 (.A ({n_514,
       n_513, n_512, n_511, n_510, n_509, n_508, n_507, n_506, n_505,
       n_504, n_503, n_502, n_501, n_500, n_499, n_498}), .B (cin), .Z
       ({n_223, n_221, n_219, n_217, n_215, n_213, n_211, n_209, n_207,
       n_205, n_203, n_201, n_199, n_197, n_195, n_193, n_191}));
  fx68k_sub_unsigned_1875 \mySubber_228_3:sub_285_24 (.A (inpb), .B
       (aOperand), .Z ({n_531, n_530, n_529, n_528, n_527, n_526,
       n_525, n_524, n_523, n_522, n_521, n_520, n_519, n_518, n_517,
       n_516, n_515}));
  fx68k_sub_signed_1877 \mySubber_228_3:sub_285_40 (.A ({n_531, n_530,
       n_529, n_528, n_527, n_526, n_525, n_524, n_523, n_522, n_521,
       n_520, n_519, n_518, n_517, n_516, n_515}), .B ({1'b0, cin}), .Z
       ({n_224, n_222, n_220, n_218, n_216, n_214, n_212, n_210, n_208,
       n_206, n_204, n_202, n_200, n_198, n_196, n_194, n_192}));
  fx68k_bmux_1882 mux_146_15(.ctl (aluAddrCtrl), .in_0 (iAddrBus),
       .in_1 (alub), .z (aOperand));
  fx68k_bmux_1883 mux_dOperand_149_9(.ctl (aluDataCtrl), .in_0
       (iDataBus), .in_1 (16'b0000000000000000), .in_2 ({_X_, _X_, _X_,
       _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_,
       _X_}), .in_3 (16'b1111111111111111), .z (inpb));
  fx68k_case_box_1144 ctl_313_16(.in_0 (oper), .out_0 ({n_153, n_154,
       n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162}));
  fx68k_mux_1884 mux_cmbsop_isShift_313_16(.ctl ({n_153, n_154, n_155,
       n_156, n_157, n_158, n_159, n_160, n_161, n_162}), .in_0
       (2'b10), .in_1 (2'b10), .in_2 (2'b11), .in_3 (2'b10), .in_4
       (2'b11), .in_5 (2'b10), .in_6 (2'b11), .in_7 (2'b10), .in_8
       (2'b11), .in_9 ({1'b0, _X_}), .z (cmbsop_isShift));
  fx68k_bmux_1882 mux_alue_433_8(.ctl (alueClkEn), .in_0
       (shftResult[31:16]), .in_1 (iDataBus), .z ({n_461, n_460, n_459,
       n_458, n_457, n_456, n_455, n_454, n_453, n_452, n_451, n_450,
       n_449, n_448, n_447, n_445}));
  fx68k_bmux_1503 mux_162_38(.ctl (isByte), .in_0 (aOperand[15]), .in_1
       (aOperand[7]), .z (n_165));
  fx68k_bmux_1503 mux_162_17(.ctl (isLong), .in_0 (n_165), .in_1
       (alue[15]), .z (shftMsb));
  fx68k_bmux_1503 mux_ccrMasked_416_14(.ctl (n_169), .in_0 (n_171),
       .in_1 (n_170), .z (ccrMasked[2]));
  fx68k_bmux_1854 mux_pswCcr_444_17(.ctl (n_167), .in_0 (ccrMasked),
       .in_1 (ftu[4:0]), .z ({n_181, n_180, n_179, n_178, n_177}));
  fx68k_bmux_1854 mux_pswCcr_442_7(.ctl (pwrUp), .in_0 ({n_181, n_180,
       n_179, n_178, n_177}), .in_1 (5'b00000), .z ({UNCONNECTED441,
       UNCONNECTED440, UNCONNECTED439, UNCONNECTED438,
       UNCONNECTED437}));
  fx68k_bmux_1503 mux_215_15(.ctl (rIrd8), .in_0 (ccr[0]), .in_1
       (n_182), .z (n_183));
  fx68k_bmux_1503 mux_shftCin_214_8(.ctl (row[7]), .in_0 (ccr[4]),
       .in_1 (n_183), .z (n_189));
  fx68k_mux_1550 mux_shftCin_205_9(.ctl ({n_184, n_185, n_186, n_187,
       n_188}), .in_0 (1'b0), .in_1 (shftMsb), .in_2 (aOperand[0]),
       .in_3 (n_189), .in_4 (aluColumn[1]), .z (shftCin));
  fx68k_bmux_1894 mux_284_13(.ctl (bAdd), .in_0 ({n_224, n_222, n_220,
       n_218, n_216, n_214, n_212, n_210, n_208, n_206, n_204, n_202,
       n_200, n_198, n_196, n_194, n_192}), .in_1 ({n_223, n_221,
       n_219, n_217, n_215, n_213, n_211, n_209, n_207, n_205, n_203,
       n_201, n_199, n_197, n_195, n_193, n_191}), .z ({n_297, n_295,
       n_293, n_291, n_289, n_287, n_285, n_283, n_281, n_279, n_277,
       n_275, n_273, n_271, n_269, n_267, n_265}));
  fx68k_bmux_1503 mux_310_18(.ctl (isByte), .in_0 (n_227), .in_1
       (n_226), .z (ccrTemp[2]));
  fx68k_bmux_1503 mux_354_20(.ctl (row[7]), .in_0 (aOperand[0]), .in_1
       (1'b0), .z (n_367));
  fx68k_bmux_1503 mux_369_30(.ctl (isByte), .in_0 (aOperand[14]), .in_1
       (aOperand[6]), .z (n_230));
  fx68k_bmux_1503 mux_369_7(.ctl (isLong), .in_0 (n_230), .in_1
       (alue[14]), .z (n_420));
  fx68k_bmux_1503 mux_292_10(.ctl (isByte), .in_0 (aOperand[15]), .in_1
       (aOperand[7]), .z (tsm));
  fx68k_bmux_1503 mux_293_10(.ctl (bAdd), .in_0 (n_231), .in_1 (tsm),
       .z (sm));
  fx68k_bmux_1503 mux_291_10(.ctl (isByte), .in_0 (inpb[15]), .in_1
       (inpb[7]), .z (dm));
  fx68k_mux_1577 mux_addCin_188_9(.ctl ({n_232, n_233, n_234, n_235}),
       .in_0 (1'b0), .in_1 (1'b1), .in_2 (ccrCore[0]), .in_3 (ccr[4]),
       .z (cin));
  fx68k_bmux_1894 mux_278_13(.ctl (bAdd), .in_0 ({n_263, n_262, n_261,
       n_260, n_259, n_258, n_257, n_255, n_253, n_251, n_249, n_247,
       n_245, n_243, n_241, n_239, n_237}), .in_1 ({6'b000000, n_256,
       n_254, n_252, n_250, n_248, n_246, n_244, n_242, n_240, n_238,
       n_236}), .z ({n_296, n_294, n_292, n_290, n_288, n_286, n_284,
       n_282, n_280, n_278, n_276, n_274, n_272, n_270, n_268, n_266,
       n_264}));
  fx68k_bmux_1894 mux_rtemp_276_8(.ctl (isByte), .in_0 ({n_297, n_295,
       n_293, n_291, n_289, n_287, n_285, n_283, n_281, n_279, n_277,
       n_275, n_273, n_271, n_269, n_267, n_265}), .in_1 ({n_296,
       n_294, n_292, n_290, n_288, n_286, n_284, n_282, n_280, n_278,
       n_276, n_274, n_272, n_270, n_268, n_266, n_264}), .z (rtemp));
  fx68k_bmux_1882 mux_result_276_8(.ctl (isByte), .in_0 ({n_295, n_293,
       n_291, n_289, n_287, n_285, n_283, n_281, n_279, n_277, n_275,
       n_273, n_271, n_269, n_267, n_265}), .in_1 ({n_278, n_278,
       n_278, n_278, n_278, n_278, n_278, n_278, n_278, n_276, n_274,
       n_272, n_270, n_268, n_266, n_264}), .z (mySubber_228_3));
  fx68k_mux_1906 mux_result_233_9(.ctl ({n_298, n_299, n_300, n_301,
       n_302, n_303, n_304}), .in_0 ({n_350, n_347, n_344, n_341,
       n_338, n_335, n_332, n_329, n_326, n_323, n_320, n_317, n_314,
       n_311, n_308, n_305}), .in_1 ({n_351, n_348, n_345, n_342,
       n_339, n_336, n_333, n_330, n_327, n_324, n_321, n_318, n_315,
       n_312, n_309, n_306}), .in_2 ({n_352, n_349, n_346, n_343,
       n_340, n_337, n_334, n_331, n_328, n_325, n_322, n_319, n_316,
       n_313, n_310, n_307}), .in_3 ({aOperand[7], aOperand[7],
       aOperand[7], aOperand[7], aOperand[7], aOperand[7], aOperand[7],
       aOperand[7], aOperand[7:0]}), .in_4 (shftResult[15:0]), .in_5
       (mySubber_228_3), .in_6 ({_X_, _X_, _X_, _X_, _X_, _X_, _X_,
       _X_, bcdLatch}), .z (result));
  fx68k_bmux_1503 mux_311_18(.ctl (isByte), .in_0 (result[15]), .in_1
       (result[7]), .z (n_353));
  fx68k_bmux_1520 mux_ccrTemp_317_18(.ctl (n_151), .in_0 ({n_353,
       1'b0}), .in_1 (2'b11), .z ({n_370, n_368}));
  fx68k_bmux_1503 mux_ccrTemp_333_26(.ctl (n_228), .in_0 (1'b0), .in_1
       (ccr[4]), .z (n_366));
  fx68k_bmux_1503 mux_cout_276_8(.ctl (isByte), .in_0 (n_297), .in_1
       (n_280), .z (subCout));
  fx68k_bmux_1503 mux_290_10(.ctl (isByte), .in_0 (n_295), .in_1
       (n_278), .z (rm));
  fx68k_mux_1926 mux_ccrTemp_313_16(.ctl ({n_354, n_355, n_356, n_357,
       n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365}), .in_0
       ({ccr[4], n_370, n_368, 1'b0}), .in_1 ({ccr[4], n_353, 2'b00}),
       .in_2 ({ccr[4], n_353, 1'b0, n_366}), .in_3 ({ccr[4], n_353,
       1'b0, aOperand[15]}), .in_4 ({shftMsb, n_353, 1'b0, shftMsb}),
       .in_5 ({aOperand[0], n_353, 1'b0, n_367}), .in_6 ({shftMsb,
       n_353, n_369, shftMsb}), .in_7 ({aOperand[0], n_353, 1'b0,
       aOperand[0]}), .in_8 ({ccr[4], n_353, 1'b0, shftMsb}), .in_9
       ({ccr[4], n_353, 1'b0, aOperand[0]}), .in_10 ({subCout, n_353,
       subOv, subCout}), .in_11 ({bcdCarry, n_353, bcdOverf,
       bcdCarry}), .z ({ccrTemp[4:3], ccrTemp[1:0]}));
  not g1 (ze, ccrCore[2]);
  not g2 (n_406, ird[6]);
  and g3 (n_407, ird[7], n_406);
  or g4 (n_408, n_407, row[7]);
  or g5 (n_411, n_408, row[1]);
  or g14 (n_404, row[7], row[1]);
  xor g18 (n_182, ccr[3], ccr[1]);
  or g19 (n_414, n_412, n_413);
  or g20 (bAdd, n_414, n_415);
  CDN_dc logicX_inst(.cf (1'b0), .dcf (1'b1), .z (_X_));
  not g25 (n_226, n_416);
  not g27 (n_227, n_417);
  or g28 (n_419, row[11], row[8]);
  xor g30 (n_421, shftMsb, n_420);
  or g31 (n_369, ccr[1], n_421);
  or g36 (n_169, finish, isArX);
  and g37 (n_170, ccrTemp[2], ccr[2]);
  and g39 (n_163, cmbsop_isShift[1], n_98);
  and g40 (n_167, enT3, ftu2Ccr);
  or g43 (n_441, finish, init);
  xor g50 (subHcarry, n_469, rtemp[4]);
  not g51 (n_471, rm);
  and g52 (n_472, n_470, n_471);
  or g53 (subOv, n_472, n_473);
  and g54 (n_473, n_474, rm);
  and g55 (n_470, sm, dm);
  not g56 (n_476, dm);
  and g57 (n_474, n_475, n_476);
  not g58 (n_475, sm);
  not g59 (n_231, tsm);
  xor g60 (n_469, aOperand[4], inpb[4]);
  not g68 (n_442, alueClkEn);
  and g79 (n_443, n_163, n_442);
  or g80 (n_444, n_443, alueClkEn);
  and g81 (n_446, n_444, enT3);
  and g82 (n_462, n_98, enT3);
  or g84 (n_465, n_464, n_167);
  CDN_flop \row_reg[0] (.clk (clk), .d (cRow[0]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[0]));
  CDN_flop \row_reg[1] (.clk (clk), .d (cRow[1]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[1]));
  CDN_flop \row_reg[2] (.clk (clk), .d (cRow[2]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[2]));
  CDN_flop \row_reg[3] (.clk (clk), .d (cRow[3]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[3]));
  CDN_flop \row_reg[4] (.clk (clk), .d (cRow[4]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[4]));
  CDN_flop \row_reg[5] (.clk (clk), .d (cRow[5]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[5]));
  CDN_flop \row_reg[6] (.clk (clk), .d (cRow[6]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[6]));
  CDN_flop \row_reg[7] (.clk (clk), .d (cRow[7]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[7]));
  CDN_flop \row_reg[8] (.clk (clk), .d (cRow[8]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[8]));
  CDN_flop \row_reg[9] (.clk (clk), .d (cRow[9]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[9]));
  CDN_flop \row_reg[10] (.clk (clk), .d (cRow[10]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[10]));
  CDN_flop \row_reg[11] (.clk (clk), .d (cRow[11]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[11]));
  CDN_flop \row_reg[12] (.clk (clk), .d (cRow[12]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[12]));
  CDN_flop \row_reg[13] (.clk (clk), .d (cRow[13]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[13]));
  CDN_flop \row_reg[14] (.clk (clk), .d (cRow[14]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[14]));
  CDN_flop \row_reg[15] (.clk (clk), .d (cRow[15]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (row[15]));
  CDN_flop isArX_reg(.clk (clk), .d (cIsArX), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (isArX));
  CDN_flop noCcrEn_reg(.clk (clk), .d (cNoCcrEn), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (noCcrEn));
  CDN_flop isByte_reg(.clk (clk), .d (aluIsByte), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (isByte));
  CDN_flop \ccrMask_reg[0] (.clk (clk), .d (cMask[0]), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ccrMask[0]));
  CDN_flop \ccrMask_reg[1] (.clk (clk), .d (cMask[1]), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ccrMask[1]));
  CDN_flop \ccrMask_reg[2] (.clk (clk), .d (cMask[2]), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ccrMask[2]));
  CDN_flop \ccrMask_reg[3] (.clk (clk), .d (cMask[3]), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ccrMask[3]));
  CDN_flop \ccrMask_reg[4] (.clk (clk), .d (cMask[4]), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ccrMask[4]));
  CDN_flop \oper_reg[0] (.clk (clk), .d (aluOp[0]), .sena (enT4), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (oper[0]));
  CDN_flop \oper_reg[1] (.clk (clk), .d (aluOp[1]), .sena (enT4), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (oper[1]));
  CDN_flop \oper_reg[2] (.clk (clk), .d (aluOp[2]), .sena (enT4), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (oper[2]));
  CDN_flop \oper_reg[3] (.clk (clk), .d (aluOp[3]), .sena (enT4), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (oper[3]));
  CDN_flop \oper_reg[4] (.clk (clk), .d (aluOp[4]), .sena (enT4), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (oper[4]));
  CDN_flop isLong_reg(.clk (clk), .d (n_411), .sena (enT4), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (isLong));
  CDN_flop rIrd8_reg(.clk (clk), .d (ird[8]), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (rIrd8));
  CDN_flop \bcdLatch_reg[0] (.clk (clk), .d (bcdResult[0]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[0]));
  CDN_flop \bcdLatch_reg[1] (.clk (clk), .d (bcdResult[1]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[1]));
  CDN_flop \bcdLatch_reg[2] (.clk (clk), .d (bcdResult[2]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[2]));
  CDN_flop \bcdLatch_reg[3] (.clk (clk), .d (bcdResult[3]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[3]));
  CDN_flop \bcdLatch_reg[4] (.clk (clk), .d (bcdResult[4]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[4]));
  CDN_flop \bcdLatch_reg[5] (.clk (clk), .d (bcdResult[5]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[5]));
  CDN_flop \bcdLatch_reg[6] (.clk (clk), .d (bcdResult[6]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[6]));
  CDN_flop \bcdLatch_reg[7] (.clk (clk), .d (bcdResult[7]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (bcdLatch[7]));
  CDN_flop bcdCarry_reg(.clk (clk), .d (bcdC), .sena (enT1), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (bcdCarry));
  CDN_flop bcdOverf_reg(.clk (clk), .d (bcdV), .sena (enT1), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (bcdOverf));
  CDN_flop \alue_reg[0] (.clk (clk), .d (n_445), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[0]));
  CDN_flop \alue_reg[1] (.clk (clk), .d (n_447), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[1]));
  CDN_flop \alue_reg[2] (.clk (clk), .d (n_448), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[2]));
  CDN_flop \alue_reg[3] (.clk (clk), .d (n_449), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[3]));
  CDN_flop \alue_reg[4] (.clk (clk), .d (n_450), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[4]));
  CDN_flop \alue_reg[5] (.clk (clk), .d (n_451), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[5]));
  CDN_flop \alue_reg[6] (.clk (clk), .d (n_452), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[6]));
  CDN_flop \alue_reg[7] (.clk (clk), .d (n_453), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[7]));
  CDN_flop \alue_reg[8] (.clk (clk), .d (n_454), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[8]));
  CDN_flop \alue_reg[9] (.clk (clk), .d (n_455), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[9]));
  CDN_flop \alue_reg[10] (.clk (clk), .d (n_456), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[10]));
  CDN_flop \alue_reg[11] (.clk (clk), .d (n_457), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[11]));
  CDN_flop \alue_reg[12] (.clk (clk), .d (n_458), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[12]));
  CDN_flop \alue_reg[13] (.clk (clk), .d (n_459), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[13]));
  CDN_flop \alue_reg[14] (.clk (clk), .d (n_460), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[14]));
  CDN_flop \alue_reg[15] (.clk (clk), .d (n_461), .sena (n_446), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (alue[15]));
  CDN_flop \aluLatch_reg[0] (.clk (clk), .d (result[0]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[0]));
  CDN_flop \aluLatch_reg[1] (.clk (clk), .d (result[1]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[1]));
  CDN_flop \aluLatch_reg[2] (.clk (clk), .d (result[2]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[2]));
  CDN_flop \aluLatch_reg[3] (.clk (clk), .d (result[3]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[3]));
  CDN_flop \aluLatch_reg[4] (.clk (clk), .d (result[4]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[4]));
  CDN_flop \aluLatch_reg[5] (.clk (clk), .d (result[5]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[5]));
  CDN_flop \aluLatch_reg[6] (.clk (clk), .d (result[6]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[6]));
  CDN_flop \aluLatch_reg[7] (.clk (clk), .d (result[7]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[7]));
  CDN_flop \aluLatch_reg[8] (.clk (clk), .d (result[8]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[8]));
  CDN_flop \aluLatch_reg[9] (.clk (clk), .d (result[9]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (aluOut[9]));
  CDN_flop \aluLatch_reg[10] (.clk (clk), .d (result[10]), .sena
       (n_462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aluOut[10]));
  CDN_flop \aluLatch_reg[11] (.clk (clk), .d (result[11]), .sena
       (n_462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aluOut[11]));
  CDN_flop \aluLatch_reg[12] (.clk (clk), .d (result[12]), .sena
       (n_462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aluOut[12]));
  CDN_flop \aluLatch_reg[13] (.clk (clk), .d (result[13]), .sena
       (n_462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aluOut[13]));
  CDN_flop \aluLatch_reg[14] (.clk (clk), .d (result[14]), .sena
       (n_462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aluOut[14]));
  CDN_flop \aluLatch_reg[15] (.clk (clk), .d (result[15]), .sena
       (n_462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aluOut[15]));
  CDN_flop \pswCcr_reg[0] (.clk (clk), .d (n_177), .sena (n_465), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ccr[0]));
  CDN_flop \pswCcr_reg[1] (.clk (clk), .d (n_178), .sena (n_465), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ccr[1]));
  CDN_flop \pswCcr_reg[2] (.clk (clk), .d (n_179), .sena (n_465), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ccr[2]));
  CDN_flop \pswCcr_reg[3] (.clk (clk), .d (n_180), .sena (n_465), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ccr[3]));
  CDN_flop \pswCcr_reg[4] (.clk (clk), .d (n_181), .sena (n_465), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ccr[4]));
  CDN_flop \ccrCore_reg[0] (.clk (clk), .d (ccrTemp[0]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ccrCore[0]));
  CDN_flop \ccrCore_reg[2] (.clk (clk), .d (ccrTemp[2]), .sena (n_462),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ccrCore[2]));
  CDN_flop coreH_reg(.clk (clk), .d (subHcarry), .sena (n_462), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (coreH));
  nand g168 (n_708, aluDataCtrl[1], n_707);
  not g169 (isCorf, n_708);
  nand g174 (n_405, n_709, oper[1], oper[2], n_712);
  nor g178 (n_712, oper[4], oper[3]);
  nand g179 (n_717, n_709, n_714, oper[2], n_712);
  not g180 (n_412, n_717);
  not g185 (n_718, oper[4]);
  nand g186 (n_723, n_718, oper[0], oper[1], n_9);
  not g187 (n_724, oper[3]);
  nor g188 (n_413, n_723, n_724);
  nand g194 (n_730, n_718, n_709, n_714, oper[2]);
  nor g196 (n_415, n_730, n_724);
  nand g200 (n_735, aluColumn[0], n_733, aluColumn[2]);
  not g201 (n_151, n_735);
  not g206 (n_709, oper[0]);
  not g207 (n_714, oper[1]);
  not g208 (n_9, oper[2]);
  not g209 (n_733, aluColumn[1]);
  not g210 (n_707, aluDataCtrl[0]);
  and g211 (n_464, n_755, n_756, enT3, n_441);
  not g212 (n_755, noCcrEn);
  not g213 (n_756, n_167);
  and g214 (n_228, n_757, n_733, aluColumn[0], n_419);
  not g215 (n_757, aluColumn[2]);
  nor g218 (n_184, n_7, n_11);
  and g220 (n_761, oper[0], oper[4]);
  and g222 (n_6, n_709, n_718);
  or g6 (n_7, n_761, n_6);
  nor g7 (n_11, n_718, n_10);
  nor g8 (n_10, oper[2], oper[1]);
  nor g9 (n_185, n_11, n_13);
  not g10 (n_13, n_7);
  nor g11 (n_186, oper[0], n_15);
  nand g12 (n_15, oper[1], oper[4]);
  nor g13 (n_187, n_17, n_21);
  not g223 (n_17, n_11);
  and g15 (n_19, oper[0], oper[2]);
  and g17 (n_20, n_709, n_9);
  or g224 (n_21, n_19, n_20);
  nor g225 (n_188, n_709, n_23);
  nand g226 (n_23, oper[2], oper[4]);
  nor g232 (n_232, oper[3], n_8);
  nand g233 (n_8, n_82, n_764);
  nand g234 (n_82, n_9, oper[0]);
  nand g236 (n_764, oper[2], oper[1]);
  not g237 (n_233, n_764);
  nor g238 (n_234, n_724, oper[2]);
  nor g240 (n_235, n_767, n_16);
  and g241 (n_766, oper[3], n_9);
  and g242 (n_14, n_724, oper[2]);
  or g243 (n_767, n_766, n_14);
  nor g244 (n_16, oper[2], oper[0]);
  nor g245 (n_298, n_775, n_777);
  nand g246 (n_775, n_718, n_724);
  nand g249 (n_777, n_714, n_9);
  nor g252 (n_299, n_12, n_779);
  nand g253 (n_12, n_718, n_9);
  nand g254 (n_779, n_714, n_709);
  nor g256 (n_300, n_780, n_781);
  nand g257 (n_780, n_714, oper[3]);
  nand g258 (n_781, oper[0], n_9);
  nor g259 (n_301, n_782, n_784);
  nand g260 (n_782, n_718, oper[2]);
  nand g261 (n_784, n_714, n_783);
  nor g262 (n_783, n_709, oper[3]);
  nor g263 (n_302, n_24, n_32);
  not g264 (n_24, n_775);
  nand g265 (n_32, n_26, n_31);
  nand g266 (n_26, n_25, n_718);
  not g267 (n_25, n_779);
  nand g268 (n_31, n_29, n_30);
  and g269 (n_27, oper[4], oper[2]);
  and g270 (n_28, n_718, n_9);
  or g271 (n_29, n_27, n_28);
  nand g272 (n_30, n_714, oper[2]);
  nor g29 (n_303, oper[4], n_42);
  nand g273 (n_42, n_39, n_786);
  nand g274 (n_39, n_37, n_38);
  nand g275 (n_37, oper[2], n_36);
  and g276 (n_34, oper[1], oper[0]);
  and g277 (n_785, n_714, n_709);
  or g278 (n_36, n_34, n_785);
  nand g279 (n_38, oper[1], n_9);
  nand g280 (n_786, oper[0], n_40);
  nor g281 (n_40, n_9, n_724);
  nor g282 (n_304, n_787, n_788);
  nand g283 (n_787, oper[1], n_724);
  nand g41 (n_788, n_709, oper[2]);
  nor g291 (n_354, n_796, n_800);
  nand g292 (n_796, n_718, oper[0]);
  nand g294 (n_800, n_724, n_799);
  nor g296 (n_799, n_9, oper[1]);
  nor g298 (n_355, n_804, n_810);
  and g299 (n_802, oper[3], oper[1]);
  and g301 (n_803, n_724, n_714);
  or g302 (n_804, n_802, n_803);
  nand g303 (n_810, n_807, n_809);
  and g304 (n_805, oper[2], oper[1]);
  and g305 (n_806, n_9, n_714);
  or g306 (n_807, n_805, n_806);
  nand g307 (n_809, n_709, oper[1]);
  nor g309 (n_356, n_811, n_812);
  nand g310 (n_811, n_718, n_714);
  nand g311 (n_812, n_724, n_9);
  nor g312 (n_357, n_718, n_813);
  nand g313 (n_813, oper[2], oper[0]);
  nor g314 (n_358, n_815, n_816);
  nor g315 (n_815, oper[4], n_814);
  nor g316 (n_814, n_724, n_9);
  nand g317 (n_816, oper[0], oper[1]);
  nor g318 (n_359, n_718, n_33);
  nand g319 (n_33, n_709, n_714);
  nor g320 (n_360, n_813, n_817);
  nand g321 (n_817, oper[3], n_714);
  nor g322 (n_361, n_818, n_819);
  nand g323 (n_818, oper[3], oper[1]);
  nand g324 (n_819, oper[2], n_709);
  nor g325 (n_362, n_820, n_82);
  nand g326 (n_820, oper[4], n_714);
  nor g328 (n_363, n_43, n_822);
  nand g329 (n_43, oper[4], oper[1]);
  nand g330 (n_822, n_9, n_709);
  nor g331 (n_364, oper[4], n_825);
  nand g332 (n_825, n_823, n_824);
  not g333 (n_823, n_807);
  nand g334 (n_824, oper[0], n_714);
  nor g335 (n_365, n_819, n_826);
  nand g336 (n_826, n_724, oper[1]);
endmodule

module fx68k_and_op_1163(A, Z);
  input [3:0] A;
  output Z;
  wire [3:0] A;
  wire Z;
  wire n_5;
  nand g1 (n_5, A[3], A[2], A[1], A[0]);
  not g2 (Z, n_5);
endmodule

module fx68k_and_op_1165(A, Z);
  input [3:0] A;
  output Z;
  wire [3:0] A;
  wire Z;
  wire n_5;
  nand g1 (n_5, A[3], A[2], A[1], A[0]);
  not g2 (Z, n_5);
endmodule

module fx68k_not_op_1232(A, Z);
  input [3:0] A;
  output [3:0] Z;
  wire [3:0] A;
  wire [3:0] Z;
  not g1 (Z[3], A[3]);
  not g2 (Z[2], A[2]);
  not g3 (Z[1], A[1]);
  not g4 (Z[0], A[0]);
endmodule

module fx68k_add_unsigned_1948(A, B, Z);
  input [31:0] A, B;
  output [31:0] Z;
  wire [31:0] A, B;
  wire [31:0] Z;
  wire n_98, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
  wire n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187;
  wire n_188, n_189, n_190, n_191, n_192, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_439;
  wire n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_98, A[0], B[0]);
  nor g6 (n_101, A[1], B[1]);
  nand g7 (n_104, A[1], B[1]);
  nor g8 (n_111, A[2], B[2]);
  nand g9 (n_106, A[2], B[2]);
  nor g10 (n_107, A[3], B[3]);
  nand g11 (n_108, A[3], B[3]);
  nor g12 (n_117, A[4], B[4]);
  nand g13 (n_112, A[4], B[4]);
  nor g14 (n_113, A[5], B[5]);
  nand g15 (n_114, A[5], B[5]);
  nor g16 (n_123, A[6], B[6]);
  nand g17 (n_118, A[6], B[6]);
  nor g18 (n_119, A[7], B[7]);
  nand g19 (n_120, A[7], B[7]);
  nor g20 (n_129, A[8], B[8]);
  nand g21 (n_124, A[8], B[8]);
  nor g22 (n_125, A[9], B[9]);
  nand g23 (n_126, A[9], B[9]);
  nor g24 (n_135, A[10], B[10]);
  nand g25 (n_130, A[10], B[10]);
  nor g26 (n_131, A[11], B[11]);
  nand g27 (n_132, A[11], B[11]);
  nor g28 (n_141, A[12], B[12]);
  nand g29 (n_136, A[12], B[12]);
  nor g30 (n_137, A[13], B[13]);
  nand g31 (n_138, A[13], B[13]);
  nor g32 (n_147, A[14], B[14]);
  nand g33 (n_142, A[14], B[14]);
  nor g34 (n_143, A[15], B[15]);
  nand g35 (n_144, A[15], B[15]);
  nor g36 (n_153, A[16], B[16]);
  nand g37 (n_148, A[16], B[16]);
  nor g38 (n_149, A[17], B[17]);
  nand g39 (n_150, A[17], B[17]);
  nor g40 (n_159, A[18], B[18]);
  nand g41 (n_154, A[18], B[18]);
  nor g42 (n_155, A[19], B[19]);
  nand g43 (n_156, A[19], B[19]);
  nor g44 (n_165, A[20], B[20]);
  nand g45 (n_160, A[20], B[20]);
  nor g46 (n_161, A[21], B[21]);
  nand g47 (n_162, A[21], B[21]);
  nor g48 (n_171, A[22], B[22]);
  nand g49 (n_166, A[22], B[22]);
  nor g50 (n_167, A[23], B[23]);
  nand g51 (n_168, A[23], B[23]);
  nor g52 (n_177, A[24], B[24]);
  nand g53 (n_172, A[24], B[24]);
  nor g54 (n_173, A[25], B[25]);
  nand g55 (n_174, A[25], B[25]);
  nor g56 (n_183, A[26], B[26]);
  nand g57 (n_178, A[26], B[26]);
  nor g58 (n_179, A[27], B[27]);
  nand g59 (n_180, A[27], B[27]);
  nor g60 (n_189, A[28], B[28]);
  nand g61 (n_184, A[28], B[28]);
  nor g62 (n_185, A[29], B[29]);
  nand g63 (n_186, A[29], B[29]);
  nor g64 (n_195, A[30], B[30]);
  nand g65 (n_190, A[30], B[30]);
  nor g66 (n_191, A[31], B[31]);
  nand g67 (n_192, A[31], B[31]);
  not g68 (n_103, n_101);
  nand g69 (n_105, n_102, n_103);
  nand g70 (n_196, n_104, n_105);
  nor g71 (n_109, n_106, n_107);
  not g72 (n_110, n_108);
  nor g73 (n_200, n_109, n_110);
  nor g74 (n_199, n_111, n_107);
  nor g75 (n_115, n_112, n_113);
  not g76 (n_116, n_114);
  nor g77 (n_202, n_115, n_116);
  nor g78 (n_205, n_117, n_113);
  nor g79 (n_121, n_118, n_119);
  not g80 (n_122, n_120);
  nor g81 (n_209, n_121, n_122);
  nor g82 (n_207, n_123, n_119);
  nor g83 (n_127, n_124, n_125);
  not g84 (n_128, n_126);
  nor g85 (n_212, n_127, n_128);
  nor g86 (n_215, n_129, n_125);
  nor g87 (n_133, n_130, n_131);
  not g88 (n_134, n_132);
  nor g89 (n_219, n_133, n_134);
  nor g90 (n_217, n_135, n_131);
  nor g91 (n_139, n_136, n_137);
  not g92 (n_140, n_138);
  nor g93 (n_222, n_139, n_140);
  nor g94 (n_225, n_141, n_137);
  nor g95 (n_145, n_142, n_143);
  not g96 (n_146, n_144);
  nor g97 (n_229, n_145, n_146);
  nor g98 (n_227, n_147, n_143);
  nor g99 (n_151, n_148, n_149);
  not g100 (n_152, n_150);
  nor g101 (n_232, n_151, n_152);
  nor g102 (n_235, n_153, n_149);
  nor g103 (n_157, n_154, n_155);
  not g104 (n_158, n_156);
  nor g105 (n_239, n_157, n_158);
  nor g106 (n_237, n_159, n_155);
  nor g107 (n_163, n_160, n_161);
  not g108 (n_164, n_162);
  nor g109 (n_242, n_163, n_164);
  nor g110 (n_245, n_165, n_161);
  nor g111 (n_169, n_166, n_167);
  not g112 (n_170, n_168);
  nor g113 (n_249, n_169, n_170);
  nor g114 (n_247, n_171, n_167);
  nor g115 (n_175, n_172, n_173);
  not g116 (n_176, n_174);
  nor g117 (n_252, n_175, n_176);
  nor g118 (n_255, n_177, n_173);
  nor g119 (n_181, n_178, n_179);
  not g120 (n_182, n_180);
  nor g121 (n_259, n_181, n_182);
  nor g122 (n_257, n_183, n_179);
  nor g123 (n_187, n_184, n_185);
  not g124 (n_188, n_186);
  nor g125 (n_262, n_187, n_188);
  nor g126 (n_265, n_189, n_185);
  not g131 (n_197, n_111);
  nand g132 (n_198, n_196, n_197);
  nand g133 (n_442, n_106, n_198);
  nand g134 (n_201, n_199, n_196);
  nand g135 (n_272, n_200, n_201);
  nor g136 (n_203, n_123, n_202);
  not g137 (n_204, n_118);
  nor g138 (n_278, n_203, n_204);
  not g139 (n_206, n_123);
  nand g140 (n_276, n_205, n_206);
  not g141 (n_208, n_207);
  nor g142 (n_210, n_202, n_208);
  not g143 (n_211, n_209);
  nor g144 (n_282, n_210, n_211);
  nand g145 (n_280, n_205, n_207);
  nor g146 (n_213, n_135, n_212);
  not g147 (n_214, n_130);
  nor g148 (n_335, n_213, n_214);
  not g149 (n_216, n_135);
  nand g150 (n_333, n_215, n_216);
  not g151 (n_218, n_217);
  nor g152 (n_220, n_212, n_218);
  not g153 (n_221, n_219);
  nor g154 (n_284, n_220, n_221);
  nand g155 (n_287, n_215, n_217);
  nor g156 (n_223, n_147, n_222);
  not g157 (n_224, n_142);
  nor g158 (n_292, n_223, n_224);
  not g159 (n_226, n_147);
  nand g160 (n_291, n_225, n_226);
  not g161 (n_228, n_227);
  nor g162 (n_230, n_222, n_228);
  not g163 (n_231, n_229);
  nor g164 (n_296, n_230, n_231);
  nand g165 (n_295, n_225, n_227);
  nor g166 (n_233, n_159, n_232);
  not g167 (n_234, n_154);
  nor g168 (n_393, n_233, n_234);
  not g169 (n_236, n_159);
  nand g170 (n_391, n_235, n_236);
  not g171 (n_238, n_237);
  nor g172 (n_240, n_232, n_238);
  not g173 (n_241, n_239);
  nor g174 (n_299, n_240, n_241);
  nand g175 (n_302, n_235, n_237);
  nor g176 (n_243, n_171, n_242);
  not g177 (n_244, n_166);
  nor g178 (n_307, n_243, n_244);
  not g179 (n_246, n_171);
  nand g180 (n_306, n_245, n_246);
  not g181 (n_248, n_247);
  nor g182 (n_250, n_242, n_248);
  not g183 (n_251, n_249);
  nor g184 (n_311, n_250, n_251);
  nand g185 (n_310, n_245, n_247);
  nor g186 (n_253, n_183, n_252);
  not g187 (n_254, n_178);
  nor g188 (n_360, n_253, n_254);
  not g189 (n_256, n_183);
  nand g190 (n_359, n_255, n_256);
  not g191 (n_258, n_257);
  nor g192 (n_260, n_252, n_258);
  not g193 (n_261, n_259);
  nor g194 (n_314, n_260, n_261);
  nand g195 (n_317, n_255, n_257);
  nor g196 (n_263, n_195, n_262);
  not g197 (n_264, n_190);
  nor g198 (n_322, n_263, n_264);
  not g199 (n_266, n_195);
  nand g200 (n_321, n_265, n_266);
  not g206 (n_273, n_117);
  nand g207 (n_274, n_272, n_273);
  nand g208 (n_446, n_112, n_274);
  nand g209 (n_275, n_205, n_272);
  nand g210 (n_448, n_202, n_275);
  not g211 (n_277, n_276);
  nand g212 (n_279, n_272, n_277);
  nand g213 (n_451, n_278, n_279);
  not g214 (n_281, n_280);
  nand g215 (n_283, n_272, n_281);
  nand g216 (n_329, n_282, n_283);
  nor g217 (n_285, n_141, n_284);
  not g218 (n_286, n_136);
  nor g219 (n_340, n_285, n_286);
  nor g220 (n_339, n_141, n_287);
  not g221 (n_288, n_225);
  nor g222 (n_289, n_284, n_288);
  not g223 (n_290, n_222);
  nor g224 (n_343, n_289, n_290);
  nor g225 (n_342, n_287, n_288);
  nor g226 (n_293, n_291, n_284);
  not g227 (n_294, n_292);
  nor g228 (n_346, n_293, n_294);
  nor g229 (n_345, n_287, n_291);
  nor g230 (n_297, n_295, n_284);
  not g231 (n_298, n_296);
  nor g232 (n_349, n_297, n_298);
  nor g233 (n_348, n_287, n_295);
  nor g234 (n_300, n_165, n_299);
  not g235 (n_301, n_160);
  nor g236 (n_398, n_300, n_301);
  nor g237 (n_397, n_165, n_302);
  not g238 (n_303, n_245);
  nor g239 (n_304, n_299, n_303);
  not g240 (n_305, n_242);
  nor g241 (n_401, n_304, n_305);
  nor g242 (n_400, n_302, n_303);
  nor g243 (n_308, n_306, n_299);
  not g244 (n_309, n_307);
  nor g245 (n_404, n_308, n_309);
  nor g246 (n_403, n_302, n_306);
  nor g247 (n_312, n_310, n_299);
  not g248 (n_313, n_311);
  nor g249 (n_351, n_312, n_313);
  nor g250 (n_354, n_302, n_310);
  nor g251 (n_315, n_189, n_314);
  not g252 (n_316, n_184);
  nor g253 (n_369, n_315, n_316);
  nor g254 (n_367, n_189, n_317);
  not g255 (n_318, n_265);
  nor g256 (n_319, n_314, n_318);
  not g257 (n_320, n_262);
  nor g258 (n_374, n_319, n_320);
  nor g259 (n_372, n_317, n_318);
  nor g260 (n_323, n_321, n_314);
  not g261 (n_324, n_322);
  nor g262 (n_379, n_323, n_324);
  nor g263 (n_377, n_317, n_321);
  not g268 (n_330, n_129);
  nand g269 (n_331, n_329, n_330);
  nand g270 (n_455, n_124, n_331);
  nand g271 (n_332, n_215, n_329);
  nand g272 (n_457, n_212, n_332);
  not g273 (n_334, n_333);
  nand g274 (n_336, n_329, n_334);
  nand g275 (n_460, n_335, n_336);
  not g276 (n_337, n_287);
  nand g277 (n_338, n_329, n_337);
  nand g278 (n_463, n_284, n_338);
  nand g279 (n_341, n_339, n_329);
  nand g280 (n_466, n_340, n_341);
  nand g281 (n_344, n_342, n_329);
  nand g282 (n_468, n_343, n_344);
  nand g283 (n_347, n_345, n_329);
  nand g284 (n_471, n_346, n_347);
  nand g285 (n_350, n_348, n_329);
  nand g286 (n_387, n_349, n_350);
  nor g287 (n_352, n_177, n_351);
  not g288 (n_353, n_172);
  nor g289 (n_409, n_352, n_353);
  not g290 (n_355, n_177);
  nand g291 (n_407, n_354, n_355);
  not g292 (n_356, n_255);
  nor g293 (n_357, n_351, n_356);
  not g294 (n_358, n_252);
  nor g295 (n_413, n_357, n_358);
  nand g296 (n_411, n_255, n_354);
  nor g297 (n_361, n_359, n_351);
  not g298 (n_362, n_360);
  nor g299 (n_417, n_361, n_362);
  not g300 (n_363, n_359);
  nand g301 (n_415, n_354, n_363);
  nor g302 (n_364, n_317, n_351);
  not g303 (n_365, n_314);
  nor g304 (n_421, n_364, n_365);
  not g305 (n_366, n_317);
  nand g306 (n_419, n_354, n_366);
  not g307 (n_368, n_367);
  nor g308 (n_370, n_351, n_368);
  not g309 (n_371, n_369);
  nor g310 (n_425, n_370, n_371);
  nand g311 (n_423, n_354, n_367);
  not g312 (n_373, n_372);
  nor g313 (n_375, n_351, n_373);
  not g314 (n_376, n_374);
  nor g315 (n_429, n_375, n_376);
  nand g316 (n_427, n_354, n_372);
  not g317 (n_378, n_377);
  nor g318 (n_380, n_351, n_378);
  not g319 (n_381, n_379);
  nor g320 (n_433, n_380, n_381);
  nand g321 (n_431, n_354, n_377);
  not g327 (n_388, n_153);
  nand g328 (n_389, n_387, n_388);
  nand g329 (n_475, n_148, n_389);
  nand g330 (n_390, n_235, n_387);
  nand g331 (n_477, n_232, n_390);
  not g332 (n_392, n_391);
  nand g333 (n_394, n_387, n_392);
  nand g334 (n_480, n_393, n_394);
  not g335 (n_395, n_302);
  nand g336 (n_396, n_387, n_395);
  nand g337 (n_483, n_299, n_396);
  nand g338 (n_399, n_397, n_387);
  nand g339 (n_486, n_398, n_399);
  nand g340 (n_402, n_400, n_387);
  nand g341 (n_488, n_401, n_402);
  nand g342 (n_405, n_403, n_387);
  nand g343 (n_491, n_404, n_405);
  nand g344 (n_406, n_354, n_387);
  nand g345 (n_493, n_351, n_406);
  not g346 (n_408, n_407);
  nand g347 (n_410, n_387, n_408);
  nand g348 (n_496, n_409, n_410);
  not g349 (n_412, n_411);
  nand g350 (n_414, n_387, n_412);
  nand g351 (n_498, n_413, n_414);
  not g352 (n_416, n_415);
  nand g353 (n_418, n_387, n_416);
  nand g354 (n_501, n_417, n_418);
  not g355 (n_420, n_419);
  nand g356 (n_422, n_387, n_420);
  nand g357 (n_504, n_421, n_422);
  not g358 (n_424, n_423);
  nand g359 (n_426, n_387, n_424);
  nand g360 (n_507, n_425, n_426);
  not g361 (n_428, n_427);
  nand g362 (n_430, n_387, n_428);
  nand g363 (n_509, n_429, n_430);
  not g364 (n_432, n_431);
  nand g365 (n_434, n_387, n_432);
  nand g366 (n_512, n_433, n_434);
  nand g370 (n_439, n_103, n_104);
  xnor g371 (Z[1], n_102, n_439);
  nand g372 (n_440, n_197, n_106);
  xnor g373 (Z[2], n_196, n_440);
  not g374 (n_441, n_107);
  nand g375 (n_443, n_441, n_108);
  xnor g376 (Z[3], n_442, n_443);
  nand g377 (n_444, n_273, n_112);
  xnor g378 (Z[4], n_272, n_444);
  not g379 (n_445, n_113);
  nand g380 (n_447, n_445, n_114);
  xnor g381 (Z[5], n_446, n_447);
  nand g382 (n_449, n_206, n_118);
  xnor g383 (Z[6], n_448, n_449);
  not g384 (n_450, n_119);
  nand g385 (n_452, n_450, n_120);
  xnor g386 (Z[7], n_451, n_452);
  nand g387 (n_453, n_330, n_124);
  xnor g388 (Z[8], n_329, n_453);
  not g389 (n_454, n_125);
  nand g390 (n_456, n_454, n_126);
  xnor g391 (Z[9], n_455, n_456);
  nand g392 (n_458, n_216, n_130);
  xnor g393 (Z[10], n_457, n_458);
  not g394 (n_459, n_131);
  nand g395 (n_461, n_459, n_132);
  xnor g396 (Z[11], n_460, n_461);
  not g397 (n_462, n_141);
  nand g398 (n_464, n_462, n_136);
  xnor g399 (Z[12], n_463, n_464);
  not g400 (n_465, n_137);
  nand g401 (n_467, n_465, n_138);
  xnor g402 (Z[13], n_466, n_467);
  nand g403 (n_469, n_226, n_142);
  xnor g404 (Z[14], n_468, n_469);
  not g405 (n_470, n_143);
  nand g406 (n_472, n_470, n_144);
  xnor g407 (Z[15], n_471, n_472);
  nand g408 (n_473, n_388, n_148);
  xnor g409 (Z[16], n_387, n_473);
  not g410 (n_474, n_149);
  nand g411 (n_476, n_474, n_150);
  xnor g412 (Z[17], n_475, n_476);
  nand g413 (n_478, n_236, n_154);
  xnor g414 (Z[18], n_477, n_478);
  not g415 (n_479, n_155);
  nand g416 (n_481, n_479, n_156);
  xnor g417 (Z[19], n_480, n_481);
  not g418 (n_482, n_165);
  nand g419 (n_484, n_482, n_160);
  xnor g420 (Z[20], n_483, n_484);
  not g421 (n_485, n_161);
  nand g422 (n_487, n_485, n_162);
  xnor g423 (Z[21], n_486, n_487);
  nand g424 (n_489, n_246, n_166);
  xnor g425 (Z[22], n_488, n_489);
  not g426 (n_490, n_167);
  nand g427 (n_492, n_490, n_168);
  xnor g428 (Z[23], n_491, n_492);
  nand g429 (n_494, n_355, n_172);
  xnor g430 (Z[24], n_493, n_494);
  not g431 (n_495, n_173);
  nand g432 (n_497, n_495, n_174);
  xnor g433 (Z[25], n_496, n_497);
  nand g434 (n_499, n_256, n_178);
  xnor g435 (Z[26], n_498, n_499);
  not g436 (n_500, n_179);
  nand g437 (n_502, n_500, n_180);
  xnor g438 (Z[27], n_501, n_502);
  not g439 (n_503, n_189);
  nand g440 (n_505, n_503, n_184);
  xnor g441 (Z[28], n_504, n_505);
  not g442 (n_506, n_185);
  nand g443 (n_508, n_506, n_186);
  xnor g444 (Z[29], n_507, n_508);
  nand g445 (n_510, n_266, n_190);
  xnor g446 (Z[30], n_509, n_510);
  not g447 (n_511, n_191);
  nand g448 (n_513, n_511, n_192);
  xnor g449 (Z[31], n_512, n_513);
  not g451 (n_102, n_98);
endmodule

module fx68k_mux_1959(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6, z);
  input [6:0] ctl;
  input in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  output z;
  wire [6:0] ctl;
  wire in_0, in_1, in_2, in_3, in_4, in_5, in_6;
  wire z;
  CDN_mux7 g1(.sel0 (ctl[6]), .data0 (in_0), .sel1 (ctl[5]), .data1
       (in_1), .sel2 (ctl[4]), .data2 (in_2), .sel3 (ctl[3]), .data3
       (in_3), .sel4 (ctl[2]), .data4 (in_4), .sel5 (ctl[1]), .data5
       (in_5), .sel6 (ctl[0]), .data6 (in_6), .z (z));
endmodule

module fx68k_bmux_1967(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16,
     in_17, z);
  input [4:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17;
  output [15:0] z;
  wire [4:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8,
       in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17;
  wire [15:0] z;
  CDN_bmux18 g1(.sel0 (ctl[0]), .data0 (in_0[15]), .data1 (in_1[15]),
       .sel1 (ctl[1]), .data2 (in_2[15]), .data3 (in_3[15]), .sel2
       (ctl[2]), .data4 (in_4[15]), .data5 (in_5[15]), .data6
       (in_6[15]), .data7 (in_7[15]), .sel3 (ctl[3]), .data8
       (in_8[15]), .data9 (in_9[15]), .data10 (in_10[15]), .data11
       (in_11[15]), .data12 (in_12[15]), .data13 (in_13[15]), .data14
       (in_14[15]), .data15 (in_15[15]), .sel4 (ctl[4]), .data16
       (in_16[15]), .data17 (in_17[15]), .z (z[15]));
  CDN_bmux18 g2(.sel0 (ctl[0]), .data0 (in_0[14]), .data1 (in_1[14]),
       .sel1 (ctl[1]), .data2 (in_2[14]), .data3 (in_3[14]), .sel2
       (ctl[2]), .data4 (in_4[14]), .data5 (in_5[14]), .data6
       (in_6[14]), .data7 (in_7[14]), .sel3 (ctl[3]), .data8
       (in_8[14]), .data9 (in_9[14]), .data10 (in_10[14]), .data11
       (in_11[14]), .data12 (in_12[14]), .data13 (in_13[14]), .data14
       (in_14[14]), .data15 (in_15[14]), .sel4 (ctl[4]), .data16
       (in_16[14]), .data17 (in_17[14]), .z (z[14]));
  CDN_bmux18 g3(.sel0 (ctl[0]), .data0 (in_0[13]), .data1 (in_1[13]),
       .sel1 (ctl[1]), .data2 (in_2[13]), .data3 (in_3[13]), .sel2
       (ctl[2]), .data4 (in_4[13]), .data5 (in_5[13]), .data6
       (in_6[13]), .data7 (in_7[13]), .sel3 (ctl[3]), .data8
       (in_8[13]), .data9 (in_9[13]), .data10 (in_10[13]), .data11
       (in_11[13]), .data12 (in_12[13]), .data13 (in_13[13]), .data14
       (in_14[13]), .data15 (in_15[13]), .sel4 (ctl[4]), .data16
       (in_16[13]), .data17 (in_17[13]), .z (z[13]));
  CDN_bmux18 g4(.sel0 (ctl[0]), .data0 (in_0[12]), .data1 (in_1[12]),
       .sel1 (ctl[1]), .data2 (in_2[12]), .data3 (in_3[12]), .sel2
       (ctl[2]), .data4 (in_4[12]), .data5 (in_5[12]), .data6
       (in_6[12]), .data7 (in_7[12]), .sel3 (ctl[3]), .data8
       (in_8[12]), .data9 (in_9[12]), .data10 (in_10[12]), .data11
       (in_11[12]), .data12 (in_12[12]), .data13 (in_13[12]), .data14
       (in_14[12]), .data15 (in_15[12]), .sel4 (ctl[4]), .data16
       (in_16[12]), .data17 (in_17[12]), .z (z[12]));
  CDN_bmux18 g5(.sel0 (ctl[0]), .data0 (in_0[11]), .data1 (in_1[11]),
       .sel1 (ctl[1]), .data2 (in_2[11]), .data3 (in_3[11]), .sel2
       (ctl[2]), .data4 (in_4[11]), .data5 (in_5[11]), .data6
       (in_6[11]), .data7 (in_7[11]), .sel3 (ctl[3]), .data8
       (in_8[11]), .data9 (in_9[11]), .data10 (in_10[11]), .data11
       (in_11[11]), .data12 (in_12[11]), .data13 (in_13[11]), .data14
       (in_14[11]), .data15 (in_15[11]), .sel4 (ctl[4]), .data16
       (in_16[11]), .data17 (in_17[11]), .z (z[11]));
  CDN_bmux18 g6(.sel0 (ctl[0]), .data0 (in_0[10]), .data1 (in_1[10]),
       .sel1 (ctl[1]), .data2 (in_2[10]), .data3 (in_3[10]), .sel2
       (ctl[2]), .data4 (in_4[10]), .data5 (in_5[10]), .data6
       (in_6[10]), .data7 (in_7[10]), .sel3 (ctl[3]), .data8
       (in_8[10]), .data9 (in_9[10]), .data10 (in_10[10]), .data11
       (in_11[10]), .data12 (in_12[10]), .data13 (in_13[10]), .data14
       (in_14[10]), .data15 (in_15[10]), .sel4 (ctl[4]), .data16
       (in_16[10]), .data17 (in_17[10]), .z (z[10]));
  CDN_bmux18 g7(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .sel2
       (ctl[2]), .data4 (in_4[9]), .data5 (in_5[9]), .data6 (in_6[9]),
       .data7 (in_7[9]), .sel3 (ctl[3]), .data8 (in_8[9]), .data9
       (in_9[9]), .data10 (in_10[9]), .data11 (in_11[9]), .data12
       (in_12[9]), .data13 (in_13[9]), .data14 (in_14[9]), .data15
       (in_15[9]), .sel4 (ctl[4]), .data16 (in_16[9]), .data17
       (in_17[9]), .z (z[9]));
  CDN_bmux18 g8(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .sel2
       (ctl[2]), .data4 (in_4[8]), .data5 (in_5[8]), .data6 (in_6[8]),
       .data7 (in_7[8]), .sel3 (ctl[3]), .data8 (in_8[8]), .data9
       (in_9[8]), .data10 (in_10[8]), .data11 (in_11[8]), .data12
       (in_12[8]), .data13 (in_13[8]), .data14 (in_14[8]), .data15
       (in_15[8]), .sel4 (ctl[4]), .data16 (in_16[8]), .data17
       (in_17[8]), .z (z[8]));
  CDN_bmux18 g9(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .data7 (in_7[7]), .sel3 (ctl[3]), .data8 (in_8[7]), .data9
       (in_9[7]), .data10 (in_10[7]), .data11 (in_11[7]), .data12
       (in_12[7]), .data13 (in_13[7]), .data14 (in_14[7]), .data15
       (in_15[7]), .sel4 (ctl[4]), .data16 (in_16[7]), .data17
       (in_17[7]), .z (z[7]));
  CDN_bmux18 g10(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .data7 (in_7[6]), .sel3 (ctl[3]), .data8 (in_8[6]), .data9
       (in_9[6]), .data10 (in_10[6]), .data11 (in_11[6]), .data12
       (in_12[6]), .data13 (in_13[6]), .data14 (in_14[6]), .data15
       (in_15[6]), .sel4 (ctl[4]), .data16 (in_16[6]), .data17
       (in_17[6]), .z (z[6]));
  CDN_bmux18 g11(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .data7 (in_7[5]), .sel3 (ctl[3]), .data8 (in_8[5]), .data9
       (in_9[5]), .data10 (in_10[5]), .data11 (in_11[5]), .data12
       (in_12[5]), .data13 (in_13[5]), .data14 (in_14[5]), .data15
       (in_15[5]), .sel4 (ctl[4]), .data16 (in_16[5]), .data17
       (in_17[5]), .z (z[5]));
  CDN_bmux18 g12(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .data7 (in_7[4]), .sel3 (ctl[3]), .data8 (in_8[4]), .data9
       (in_9[4]), .data10 (in_10[4]), .data11 (in_11[4]), .data12
       (in_12[4]), .data13 (in_13[4]), .data14 (in_14[4]), .data15
       (in_15[4]), .sel4 (ctl[4]), .data16 (in_16[4]), .data17
       (in_17[4]), .z (z[4]));
  CDN_bmux18 g13(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .sel3 (ctl[3]), .data8 (in_8[3]), .data9
       (in_9[3]), .data10 (in_10[3]), .data11 (in_11[3]), .data12
       (in_12[3]), .data13 (in_13[3]), .data14 (in_14[3]), .data15
       (in_15[3]), .sel4 (ctl[4]), .data16 (in_16[3]), .data17
       (in_17[3]), .z (z[3]));
  CDN_bmux18 g14(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .sel3 (ctl[3]), .data8 (in_8[2]), .data9
       (in_9[2]), .data10 (in_10[2]), .data11 (in_11[2]), .data12
       (in_12[2]), .data13 (in_13[2]), .data14 (in_14[2]), .data15
       (in_15[2]), .sel4 (ctl[4]), .data16 (in_16[2]), .data17
       (in_17[2]), .z (z[2]));
  CDN_bmux18 g15(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .sel3 (ctl[3]), .data8 (in_8[1]), .data9
       (in_9[1]), .data10 (in_10[1]), .data11 (in_11[1]), .data12
       (in_12[1]), .data13 (in_13[1]), .data14 (in_14[1]), .data15
       (in_15[1]), .sel4 (ctl[4]), .data16 (in_16[1]), .data17
       (in_17[1]), .z (z[1]));
  CDN_bmux18 g16(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .sel3 (ctl[3]), .data8 (in_8[0]), .data9
       (in_9[0]), .data10 (in_10[0]), .data11 (in_11[0]), .data12
       (in_12[0]), .data13 (in_13[0]), .data14 (in_14[0]), .data15
       (in_15[0]), .sel4 (ctl[4]), .data16 (in_16[0]), .data17
       (in_17[0]), .z (z[0]));
endmodule

module fx68k_mux_1995(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input [15:0] in_0, in_1;
  output [15:0] z;
  wire [1:0] ctl;
  wire [15:0] in_0, in_1;
  wire [15:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[15]), .sel1 (ctl[0]), .data1
       (in_1[15]), .z (z[15]));
  CDN_mux2 g17(.sel0 (ctl[1]), .data0 (in_0[14]), .sel1 (ctl[0]),
       .data1 (in_1[14]), .z (z[14]));
  CDN_mux2 g18(.sel0 (ctl[1]), .data0 (in_0[13]), .sel1 (ctl[0]),
       .data1 (in_1[13]), .z (z[13]));
  CDN_mux2 g19(.sel0 (ctl[1]), .data0 (in_0[12]), .sel1 (ctl[0]),
       .data1 (in_1[12]), .z (z[12]));
  CDN_mux2 g20(.sel0 (ctl[1]), .data0 (in_0[11]), .sel1 (ctl[0]),
       .data1 (in_1[11]), .z (z[11]));
  CDN_mux2 g21(.sel0 (ctl[1]), .data0 (in_0[10]), .sel1 (ctl[0]),
       .data1 (in_1[10]), .z (z[10]));
  CDN_mux2 g22(.sel0 (ctl[1]), .data0 (in_0[9]), .sel1 (ctl[0]), .data1
       (in_1[9]), .z (z[9]));
  CDN_mux2 g23(.sel0 (ctl[1]), .data0 (in_0[8]), .sel1 (ctl[0]), .data1
       (in_1[8]), .z (z[8]));
  CDN_mux2 g24(.sel0 (ctl[1]), .data0 (in_0[7]), .sel1 (ctl[0]), .data1
       (in_1[7]), .z (z[7]));
  CDN_mux2 g25(.sel0 (ctl[1]), .data0 (in_0[6]), .sel1 (ctl[0]), .data1
       (in_1[6]), .z (z[6]));
  CDN_mux2 g26(.sel0 (ctl[1]), .data0 (in_0[5]), .sel1 (ctl[0]), .data1
       (in_1[5]), .z (z[5]));
  CDN_mux2 g27(.sel0 (ctl[1]), .data0 (in_0[4]), .sel1 (ctl[0]), .data1
       (in_1[4]), .z (z[4]));
  CDN_mux2 g28(.sel0 (ctl[1]), .data0 (in_0[3]), .sel1 (ctl[0]), .data1
       (in_1[3]), .z (z[3]));
  CDN_mux2 g29(.sel0 (ctl[1]), .data0 (in_0[2]), .sel1 (ctl[0]), .data1
       (in_1[2]), .z (z[2]));
  CDN_mux2 g30(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g31(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_mux_2286(ctl, in_0, in_1, in_2, in_3, in_4, z);
  input [4:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3, in_4;
  output [15:0] z;
  wire [4:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3, in_4;
  wire [15:0] z;
  CDN_mux5 g1(.sel0 (ctl[4]), .data0 (in_0[15]), .sel1 (ctl[3]), .data1
       (in_1[15]), .sel2 (ctl[2]), .data2 (in_2[15]), .sel3 (ctl[1]),
       .data3 (in_3[15]), .sel4 (ctl[0]), .data4 (in_4[15]), .z
       (z[15]));
  CDN_mux5 g17(.sel0 (ctl[4]), .data0 (in_0[14]), .sel1 (ctl[3]),
       .data1 (in_1[14]), .sel2 (ctl[2]), .data2 (in_2[14]), .sel3
       (ctl[1]), .data3 (in_3[14]), .sel4 (ctl[0]), .data4 (in_4[14]),
       .z (z[14]));
  CDN_mux5 g18(.sel0 (ctl[4]), .data0 (in_0[13]), .sel1 (ctl[3]),
       .data1 (in_1[13]), .sel2 (ctl[2]), .data2 (in_2[13]), .sel3
       (ctl[1]), .data3 (in_3[13]), .sel4 (ctl[0]), .data4 (in_4[13]),
       .z (z[13]));
  CDN_mux5 g19(.sel0 (ctl[4]), .data0 (in_0[12]), .sel1 (ctl[3]),
       .data1 (in_1[12]), .sel2 (ctl[2]), .data2 (in_2[12]), .sel3
       (ctl[1]), .data3 (in_3[12]), .sel4 (ctl[0]), .data4 (in_4[12]),
       .z (z[12]));
  CDN_mux5 g20(.sel0 (ctl[4]), .data0 (in_0[11]), .sel1 (ctl[3]),
       .data1 (in_1[11]), .sel2 (ctl[2]), .data2 (in_2[11]), .sel3
       (ctl[1]), .data3 (in_3[11]), .sel4 (ctl[0]), .data4 (in_4[11]),
       .z (z[11]));
  CDN_mux5 g21(.sel0 (ctl[4]), .data0 (in_0[10]), .sel1 (ctl[3]),
       .data1 (in_1[10]), .sel2 (ctl[2]), .data2 (in_2[10]), .sel3
       (ctl[1]), .data3 (in_3[10]), .sel4 (ctl[0]), .data4 (in_4[10]),
       .z (z[10]));
  CDN_mux5 g22(.sel0 (ctl[4]), .data0 (in_0[9]), .sel1 (ctl[3]), .data1
       (in_1[9]), .sel2 (ctl[2]), .data2 (in_2[9]), .sel3 (ctl[1]),
       .data3 (in_3[9]), .sel4 (ctl[0]), .data4 (in_4[9]), .z (z[9]));
  CDN_mux5 g23(.sel0 (ctl[4]), .data0 (in_0[8]), .sel1 (ctl[3]), .data1
       (in_1[8]), .sel2 (ctl[2]), .data2 (in_2[8]), .sel3 (ctl[1]),
       .data3 (in_3[8]), .sel4 (ctl[0]), .data4 (in_4[8]), .z (z[8]));
  CDN_mux5 g24(.sel0 (ctl[4]), .data0 (in_0[7]), .sel1 (ctl[3]), .data1
       (in_1[7]), .sel2 (ctl[2]), .data2 (in_2[7]), .sel3 (ctl[1]),
       .data3 (in_3[7]), .sel4 (ctl[0]), .data4 (in_4[7]), .z (z[7]));
  CDN_mux5 g25(.sel0 (ctl[4]), .data0 (in_0[6]), .sel1 (ctl[3]), .data1
       (in_1[6]), .sel2 (ctl[2]), .data2 (in_2[6]), .sel3 (ctl[1]),
       .data3 (in_3[6]), .sel4 (ctl[0]), .data4 (in_4[6]), .z (z[6]));
  CDN_mux5 g26(.sel0 (ctl[4]), .data0 (in_0[5]), .sel1 (ctl[3]), .data1
       (in_1[5]), .sel2 (ctl[2]), .data2 (in_2[5]), .sel3 (ctl[1]),
       .data3 (in_3[5]), .sel4 (ctl[0]), .data4 (in_4[5]), .z (z[5]));
  CDN_mux5 g27(.sel0 (ctl[4]), .data0 (in_0[4]), .sel1 (ctl[3]), .data1
       (in_1[4]), .sel2 (ctl[2]), .data2 (in_2[4]), .sel3 (ctl[1]),
       .data3 (in_3[4]), .sel4 (ctl[0]), .data4 (in_4[4]), .z (z[4]));
  CDN_mux5 g28(.sel0 (ctl[4]), .data0 (in_0[3]), .sel1 (ctl[3]), .data1
       (in_1[3]), .sel2 (ctl[2]), .data2 (in_2[3]), .sel3 (ctl[1]),
       .data3 (in_3[3]), .sel4 (ctl[0]), .data4 (in_4[3]), .z (z[3]));
  CDN_mux5 g29(.sel0 (ctl[4]), .data0 (in_0[2]), .sel1 (ctl[3]), .data1
       (in_1[2]), .sel2 (ctl[2]), .data2 (in_2[2]), .sel3 (ctl[1]),
       .data3 (in_3[2]), .sel4 (ctl[0]), .data4 (in_4[2]), .z (z[2]));
  CDN_mux5 g30(.sel0 (ctl[4]), .data0 (in_0[1]), .sel1 (ctl[3]), .data1
       (in_1[1]), .sel2 (ctl[2]), .data2 (in_2[1]), .sel3 (ctl[1]),
       .data3 (in_3[1]), .sel4 (ctl[0]), .data4 (in_4[1]), .z (z[1]));
  CDN_mux5 g31(.sel0 (ctl[4]), .data0 (in_0[0]), .sel1 (ctl[3]), .data1
       (in_1[0]), .sel2 (ctl[2]), .data2 (in_2[0]), .sel3 (ctl[1]),
       .data3 (in_3[0]), .sel4 (ctl[0]), .data4 (in_4[0]), .z (z[0]));
endmodule

module fx68k_mux_2306(ctl, in_0, in_1, in_2, in_3, in_4, in_5, z);
  input [5:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3, in_4, in_5;
  output [15:0] z;
  wire [5:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3, in_4, in_5;
  wire [15:0] z;
  CDN_mux6 g1(.sel0 (ctl[5]), .data0 (in_0[15]), .sel1 (ctl[4]), .data1
       (in_1[15]), .sel2 (ctl[3]), .data2 (in_2[15]), .sel3 (ctl[2]),
       .data3 (in_3[15]), .sel4 (ctl[1]), .data4 (in_4[15]), .sel5
       (ctl[0]), .data5 (in_5[15]), .z (z[15]));
  CDN_mux6 g17(.sel0 (ctl[5]), .data0 (in_0[14]), .sel1 (ctl[4]),
       .data1 (in_1[14]), .sel2 (ctl[3]), .data2 (in_2[14]), .sel3
       (ctl[2]), .data3 (in_3[14]), .sel4 (ctl[1]), .data4 (in_4[14]),
       .sel5 (ctl[0]), .data5 (in_5[14]), .z (z[14]));
  CDN_mux6 g18(.sel0 (ctl[5]), .data0 (in_0[13]), .sel1 (ctl[4]),
       .data1 (in_1[13]), .sel2 (ctl[3]), .data2 (in_2[13]), .sel3
       (ctl[2]), .data3 (in_3[13]), .sel4 (ctl[1]), .data4 (in_4[13]),
       .sel5 (ctl[0]), .data5 (in_5[13]), .z (z[13]));
  CDN_mux6 g19(.sel0 (ctl[5]), .data0 (in_0[12]), .sel1 (ctl[4]),
       .data1 (in_1[12]), .sel2 (ctl[3]), .data2 (in_2[12]), .sel3
       (ctl[2]), .data3 (in_3[12]), .sel4 (ctl[1]), .data4 (in_4[12]),
       .sel5 (ctl[0]), .data5 (in_5[12]), .z (z[12]));
  CDN_mux6 g20(.sel0 (ctl[5]), .data0 (in_0[11]), .sel1 (ctl[4]),
       .data1 (in_1[11]), .sel2 (ctl[3]), .data2 (in_2[11]), .sel3
       (ctl[2]), .data3 (in_3[11]), .sel4 (ctl[1]), .data4 (in_4[11]),
       .sel5 (ctl[0]), .data5 (in_5[11]), .z (z[11]));
  CDN_mux6 g21(.sel0 (ctl[5]), .data0 (in_0[10]), .sel1 (ctl[4]),
       .data1 (in_1[10]), .sel2 (ctl[3]), .data2 (in_2[10]), .sel3
       (ctl[2]), .data3 (in_3[10]), .sel4 (ctl[1]), .data4 (in_4[10]),
       .sel5 (ctl[0]), .data5 (in_5[10]), .z (z[10]));
  CDN_mux6 g22(.sel0 (ctl[5]), .data0 (in_0[9]), .sel1 (ctl[4]), .data1
       (in_1[9]), .sel2 (ctl[3]), .data2 (in_2[9]), .sel3 (ctl[2]),
       .data3 (in_3[9]), .sel4 (ctl[1]), .data4 (in_4[9]), .sel5
       (ctl[0]), .data5 (in_5[9]), .z (z[9]));
  CDN_mux6 g23(.sel0 (ctl[5]), .data0 (in_0[8]), .sel1 (ctl[4]), .data1
       (in_1[8]), .sel2 (ctl[3]), .data2 (in_2[8]), .sel3 (ctl[2]),
       .data3 (in_3[8]), .sel4 (ctl[1]), .data4 (in_4[8]), .sel5
       (ctl[0]), .data5 (in_5[8]), .z (z[8]));
  CDN_mux6 g24(.sel0 (ctl[5]), .data0 (in_0[7]), .sel1 (ctl[4]), .data1
       (in_1[7]), .sel2 (ctl[3]), .data2 (in_2[7]), .sel3 (ctl[2]),
       .data3 (in_3[7]), .sel4 (ctl[1]), .data4 (in_4[7]), .sel5
       (ctl[0]), .data5 (in_5[7]), .z (z[7]));
  CDN_mux6 g25(.sel0 (ctl[5]), .data0 (in_0[6]), .sel1 (ctl[4]), .data1
       (in_1[6]), .sel2 (ctl[3]), .data2 (in_2[6]), .sel3 (ctl[2]),
       .data3 (in_3[6]), .sel4 (ctl[1]), .data4 (in_4[6]), .sel5
       (ctl[0]), .data5 (in_5[6]), .z (z[6]));
  CDN_mux6 g26(.sel0 (ctl[5]), .data0 (in_0[5]), .sel1 (ctl[4]), .data1
       (in_1[5]), .sel2 (ctl[3]), .data2 (in_2[5]), .sel3 (ctl[2]),
       .data3 (in_3[5]), .sel4 (ctl[1]), .data4 (in_4[5]), .sel5
       (ctl[0]), .data5 (in_5[5]), .z (z[5]));
  CDN_mux6 g27(.sel0 (ctl[5]), .data0 (in_0[4]), .sel1 (ctl[4]), .data1
       (in_1[4]), .sel2 (ctl[3]), .data2 (in_2[4]), .sel3 (ctl[2]),
       .data3 (in_3[4]), .sel4 (ctl[1]), .data4 (in_4[4]), .sel5
       (ctl[0]), .data5 (in_5[4]), .z (z[4]));
  CDN_mux6 g28(.sel0 (ctl[5]), .data0 (in_0[3]), .sel1 (ctl[4]), .data1
       (in_1[3]), .sel2 (ctl[3]), .data2 (in_2[3]), .sel3 (ctl[2]),
       .data3 (in_3[3]), .sel4 (ctl[1]), .data4 (in_4[3]), .sel5
       (ctl[0]), .data5 (in_5[3]), .z (z[3]));
  CDN_mux6 g29(.sel0 (ctl[5]), .data0 (in_0[2]), .sel1 (ctl[4]), .data1
       (in_1[2]), .sel2 (ctl[3]), .data2 (in_2[2]), .sel3 (ctl[2]),
       .data3 (in_3[2]), .sel4 (ctl[1]), .data4 (in_4[2]), .sel5
       (ctl[0]), .data5 (in_5[2]), .z (z[2]));
  CDN_mux6 g30(.sel0 (ctl[5]), .data0 (in_0[1]), .sel1 (ctl[4]), .data1
       (in_1[1]), .sel2 (ctl[3]), .data2 (in_2[1]), .sel3 (ctl[2]),
       .data3 (in_3[1]), .sel4 (ctl[1]), .data4 (in_4[1]), .sel5
       (ctl[0]), .data5 (in_5[1]), .z (z[1]));
  CDN_mux6 g31(.sel0 (ctl[5]), .data0 (in_0[0]), .sel1 (ctl[4]), .data1
       (in_1[0]), .sel2 (ctl[3]), .data2 (in_2[0]), .sel3 (ctl[2]),
       .data3 (in_3[0]), .sel4 (ctl[1]), .data4 (in_4[0]), .sel5
       (ctl[0]), .data5 (in_5[0]), .z (z[0]));
endmodule

module fx68k_mux_2324(ctl, in_0, in_1, in_2, in_3, z);
  input [3:0] ctl;
  input [15:0] in_0, in_1, in_2, in_3;
  output [15:0] z;
  wire [3:0] ctl;
  wire [15:0] in_0, in_1, in_2, in_3;
  wire [15:0] z;
  CDN_mux4 g1(.sel0 (ctl[3]), .data0 (in_0[15]), .sel1 (ctl[2]), .data1
       (in_1[15]), .sel2 (ctl[1]), .data2 (in_2[15]), .sel3 (ctl[0]),
       .data3 (in_3[15]), .z (z[15]));
  CDN_mux4 g17(.sel0 (ctl[3]), .data0 (in_0[14]), .sel1 (ctl[2]),
       .data1 (in_1[14]), .sel2 (ctl[1]), .data2 (in_2[14]), .sel3
       (ctl[0]), .data3 (in_3[14]), .z (z[14]));
  CDN_mux4 g18(.sel0 (ctl[3]), .data0 (in_0[13]), .sel1 (ctl[2]),
       .data1 (in_1[13]), .sel2 (ctl[1]), .data2 (in_2[13]), .sel3
       (ctl[0]), .data3 (in_3[13]), .z (z[13]));
  CDN_mux4 g19(.sel0 (ctl[3]), .data0 (in_0[12]), .sel1 (ctl[2]),
       .data1 (in_1[12]), .sel2 (ctl[1]), .data2 (in_2[12]), .sel3
       (ctl[0]), .data3 (in_3[12]), .z (z[12]));
  CDN_mux4 g20(.sel0 (ctl[3]), .data0 (in_0[11]), .sel1 (ctl[2]),
       .data1 (in_1[11]), .sel2 (ctl[1]), .data2 (in_2[11]), .sel3
       (ctl[0]), .data3 (in_3[11]), .z (z[11]));
  CDN_mux4 g21(.sel0 (ctl[3]), .data0 (in_0[10]), .sel1 (ctl[2]),
       .data1 (in_1[10]), .sel2 (ctl[1]), .data2 (in_2[10]), .sel3
       (ctl[0]), .data3 (in_3[10]), .z (z[10]));
  CDN_mux4 g22(.sel0 (ctl[3]), .data0 (in_0[9]), .sel1 (ctl[2]), .data1
       (in_1[9]), .sel2 (ctl[1]), .data2 (in_2[9]), .sel3 (ctl[0]),
       .data3 (in_3[9]), .z (z[9]));
  CDN_mux4 g23(.sel0 (ctl[3]), .data0 (in_0[8]), .sel1 (ctl[2]), .data1
       (in_1[8]), .sel2 (ctl[1]), .data2 (in_2[8]), .sel3 (ctl[0]),
       .data3 (in_3[8]), .z (z[8]));
  CDN_mux4 g24(.sel0 (ctl[3]), .data0 (in_0[7]), .sel1 (ctl[2]), .data1
       (in_1[7]), .sel2 (ctl[1]), .data2 (in_2[7]), .sel3 (ctl[0]),
       .data3 (in_3[7]), .z (z[7]));
  CDN_mux4 g25(.sel0 (ctl[3]), .data0 (in_0[6]), .sel1 (ctl[2]), .data1
       (in_1[6]), .sel2 (ctl[1]), .data2 (in_2[6]), .sel3 (ctl[0]),
       .data3 (in_3[6]), .z (z[6]));
  CDN_mux4 g26(.sel0 (ctl[3]), .data0 (in_0[5]), .sel1 (ctl[2]), .data1
       (in_1[5]), .sel2 (ctl[1]), .data2 (in_2[5]), .sel3 (ctl[0]),
       .data3 (in_3[5]), .z (z[5]));
  CDN_mux4 g27(.sel0 (ctl[3]), .data0 (in_0[4]), .sel1 (ctl[2]), .data1
       (in_1[4]), .sel2 (ctl[1]), .data2 (in_2[4]), .sel3 (ctl[0]),
       .data3 (in_3[4]), .z (z[4]));
  CDN_mux4 g28(.sel0 (ctl[3]), .data0 (in_0[3]), .sel1 (ctl[2]), .data1
       (in_1[3]), .sel2 (ctl[1]), .data2 (in_2[3]), .sel3 (ctl[0]),
       .data3 (in_3[3]), .z (z[3]));
  CDN_mux4 g29(.sel0 (ctl[3]), .data0 (in_0[2]), .sel1 (ctl[2]), .data1
       (in_1[2]), .sel2 (ctl[1]), .data2 (in_2[2]), .sel3 (ctl[0]),
       .data3 (in_3[2]), .z (z[2]));
  CDN_mux4 g30(.sel0 (ctl[3]), .data0 (in_0[1]), .sel1 (ctl[2]), .data1
       (in_1[1]), .sel2 (ctl[1]), .data2 (in_2[1]), .sel3 (ctl[0]),
       .data3 (in_3[1]), .z (z[1]));
  CDN_mux4 g31(.sel0 (ctl[3]), .data0 (in_0[0]), .sel1 (ctl[2]), .data1
       (in_1[0]), .sel2 (ctl[1]), .data2 (in_2[0]), .sel3 (ctl[0]),
       .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_bmux_2394(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, z);
  input [2:0] ctl;
  input [31:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  output [31:0] z;
  wire [2:0] ctl;
  wire [31:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
  wire [31:0] z;
  CDN_bmux8 g1(.sel0 (ctl[0]), .data0 (in_0[31]), .data1 (in_1[31]),
       .sel1 (ctl[1]), .data2 (in_2[31]), .data3 (in_3[31]), .sel2
       (ctl[2]), .data4 (in_4[31]), .data5 (in_5[31]), .data6
       (in_6[31]), .data7 (in_7[31]), .z (z[31]));
  CDN_bmux8 g2(.sel0 (ctl[0]), .data0 (in_0[30]), .data1 (in_1[30]),
       .sel1 (ctl[1]), .data2 (in_2[30]), .data3 (in_3[30]), .sel2
       (ctl[2]), .data4 (in_4[30]), .data5 (in_5[30]), .data6
       (in_6[30]), .data7 (in_7[30]), .z (z[30]));
  CDN_bmux8 g3(.sel0 (ctl[0]), .data0 (in_0[29]), .data1 (in_1[29]),
       .sel1 (ctl[1]), .data2 (in_2[29]), .data3 (in_3[29]), .sel2
       (ctl[2]), .data4 (in_4[29]), .data5 (in_5[29]), .data6
       (in_6[29]), .data7 (in_7[29]), .z (z[29]));
  CDN_bmux8 g4(.sel0 (ctl[0]), .data0 (in_0[28]), .data1 (in_1[28]),
       .sel1 (ctl[1]), .data2 (in_2[28]), .data3 (in_3[28]), .sel2
       (ctl[2]), .data4 (in_4[28]), .data5 (in_5[28]), .data6
       (in_6[28]), .data7 (in_7[28]), .z (z[28]));
  CDN_bmux8 g5(.sel0 (ctl[0]), .data0 (in_0[27]), .data1 (in_1[27]),
       .sel1 (ctl[1]), .data2 (in_2[27]), .data3 (in_3[27]), .sel2
       (ctl[2]), .data4 (in_4[27]), .data5 (in_5[27]), .data6
       (in_6[27]), .data7 (in_7[27]), .z (z[27]));
  CDN_bmux8 g6(.sel0 (ctl[0]), .data0 (in_0[26]), .data1 (in_1[26]),
       .sel1 (ctl[1]), .data2 (in_2[26]), .data3 (in_3[26]), .sel2
       (ctl[2]), .data4 (in_4[26]), .data5 (in_5[26]), .data6
       (in_6[26]), .data7 (in_7[26]), .z (z[26]));
  CDN_bmux8 g7(.sel0 (ctl[0]), .data0 (in_0[25]), .data1 (in_1[25]),
       .sel1 (ctl[1]), .data2 (in_2[25]), .data3 (in_3[25]), .sel2
       (ctl[2]), .data4 (in_4[25]), .data5 (in_5[25]), .data6
       (in_6[25]), .data7 (in_7[25]), .z (z[25]));
  CDN_bmux8 g8(.sel0 (ctl[0]), .data0 (in_0[24]), .data1 (in_1[24]),
       .sel1 (ctl[1]), .data2 (in_2[24]), .data3 (in_3[24]), .sel2
       (ctl[2]), .data4 (in_4[24]), .data5 (in_5[24]), .data6
       (in_6[24]), .data7 (in_7[24]), .z (z[24]));
  CDN_bmux8 g9(.sel0 (ctl[0]), .data0 (in_0[23]), .data1 (in_1[23]),
       .sel1 (ctl[1]), .data2 (in_2[23]), .data3 (in_3[23]), .sel2
       (ctl[2]), .data4 (in_4[23]), .data5 (in_5[23]), .data6
       (in_6[23]), .data7 (in_7[23]), .z (z[23]));
  CDN_bmux8 g10(.sel0 (ctl[0]), .data0 (in_0[22]), .data1 (in_1[22]),
       .sel1 (ctl[1]), .data2 (in_2[22]), .data3 (in_3[22]), .sel2
       (ctl[2]), .data4 (in_4[22]), .data5 (in_5[22]), .data6
       (in_6[22]), .data7 (in_7[22]), .z (z[22]));
  CDN_bmux8 g11(.sel0 (ctl[0]), .data0 (in_0[21]), .data1 (in_1[21]),
       .sel1 (ctl[1]), .data2 (in_2[21]), .data3 (in_3[21]), .sel2
       (ctl[2]), .data4 (in_4[21]), .data5 (in_5[21]), .data6
       (in_6[21]), .data7 (in_7[21]), .z (z[21]));
  CDN_bmux8 g12(.sel0 (ctl[0]), .data0 (in_0[20]), .data1 (in_1[20]),
       .sel1 (ctl[1]), .data2 (in_2[20]), .data3 (in_3[20]), .sel2
       (ctl[2]), .data4 (in_4[20]), .data5 (in_5[20]), .data6
       (in_6[20]), .data7 (in_7[20]), .z (z[20]));
  CDN_bmux8 g13(.sel0 (ctl[0]), .data0 (in_0[19]), .data1 (in_1[19]),
       .sel1 (ctl[1]), .data2 (in_2[19]), .data3 (in_3[19]), .sel2
       (ctl[2]), .data4 (in_4[19]), .data5 (in_5[19]), .data6
       (in_6[19]), .data7 (in_7[19]), .z (z[19]));
  CDN_bmux8 g14(.sel0 (ctl[0]), .data0 (in_0[18]), .data1 (in_1[18]),
       .sel1 (ctl[1]), .data2 (in_2[18]), .data3 (in_3[18]), .sel2
       (ctl[2]), .data4 (in_4[18]), .data5 (in_5[18]), .data6
       (in_6[18]), .data7 (in_7[18]), .z (z[18]));
  CDN_bmux8 g15(.sel0 (ctl[0]), .data0 (in_0[17]), .data1 (in_1[17]),
       .sel1 (ctl[1]), .data2 (in_2[17]), .data3 (in_3[17]), .sel2
       (ctl[2]), .data4 (in_4[17]), .data5 (in_5[17]), .data6
       (in_6[17]), .data7 (in_7[17]), .z (z[17]));
  CDN_bmux8 g16(.sel0 (ctl[0]), .data0 (in_0[16]), .data1 (in_1[16]),
       .sel1 (ctl[1]), .data2 (in_2[16]), .data3 (in_3[16]), .sel2
       (ctl[2]), .data4 (in_4[16]), .data5 (in_5[16]), .data6
       (in_6[16]), .data7 (in_7[16]), .z (z[16]));
  CDN_bmux8 g17(.sel0 (ctl[0]), .data0 (in_0[15]), .data1 (in_1[15]),
       .sel1 (ctl[1]), .data2 (in_2[15]), .data3 (in_3[15]), .sel2
       (ctl[2]), .data4 (in_4[15]), .data5 (in_5[15]), .data6
       (in_6[15]), .data7 (in_7[15]), .z (z[15]));
  CDN_bmux8 g18(.sel0 (ctl[0]), .data0 (in_0[14]), .data1 (in_1[14]),
       .sel1 (ctl[1]), .data2 (in_2[14]), .data3 (in_3[14]), .sel2
       (ctl[2]), .data4 (in_4[14]), .data5 (in_5[14]), .data6
       (in_6[14]), .data7 (in_7[14]), .z (z[14]));
  CDN_bmux8 g19(.sel0 (ctl[0]), .data0 (in_0[13]), .data1 (in_1[13]),
       .sel1 (ctl[1]), .data2 (in_2[13]), .data3 (in_3[13]), .sel2
       (ctl[2]), .data4 (in_4[13]), .data5 (in_5[13]), .data6
       (in_6[13]), .data7 (in_7[13]), .z (z[13]));
  CDN_bmux8 g20(.sel0 (ctl[0]), .data0 (in_0[12]), .data1 (in_1[12]),
       .sel1 (ctl[1]), .data2 (in_2[12]), .data3 (in_3[12]), .sel2
       (ctl[2]), .data4 (in_4[12]), .data5 (in_5[12]), .data6
       (in_6[12]), .data7 (in_7[12]), .z (z[12]));
  CDN_bmux8 g21(.sel0 (ctl[0]), .data0 (in_0[11]), .data1 (in_1[11]),
       .sel1 (ctl[1]), .data2 (in_2[11]), .data3 (in_3[11]), .sel2
       (ctl[2]), .data4 (in_4[11]), .data5 (in_5[11]), .data6
       (in_6[11]), .data7 (in_7[11]), .z (z[11]));
  CDN_bmux8 g22(.sel0 (ctl[0]), .data0 (in_0[10]), .data1 (in_1[10]),
       .sel1 (ctl[1]), .data2 (in_2[10]), .data3 (in_3[10]), .sel2
       (ctl[2]), .data4 (in_4[10]), .data5 (in_5[10]), .data6
       (in_6[10]), .data7 (in_7[10]), .z (z[10]));
  CDN_bmux8 g23(.sel0 (ctl[0]), .data0 (in_0[9]), .data1 (in_1[9]),
       .sel1 (ctl[1]), .data2 (in_2[9]), .data3 (in_3[9]), .sel2
       (ctl[2]), .data4 (in_4[9]), .data5 (in_5[9]), .data6 (in_6[9]),
       .data7 (in_7[9]), .z (z[9]));
  CDN_bmux8 g24(.sel0 (ctl[0]), .data0 (in_0[8]), .data1 (in_1[8]),
       .sel1 (ctl[1]), .data2 (in_2[8]), .data3 (in_3[8]), .sel2
       (ctl[2]), .data4 (in_4[8]), .data5 (in_5[8]), .data6 (in_6[8]),
       .data7 (in_7[8]), .z (z[8]));
  CDN_bmux8 g25(.sel0 (ctl[0]), .data0 (in_0[7]), .data1 (in_1[7]),
       .sel1 (ctl[1]), .data2 (in_2[7]), .data3 (in_3[7]), .sel2
       (ctl[2]), .data4 (in_4[7]), .data5 (in_5[7]), .data6 (in_6[7]),
       .data7 (in_7[7]), .z (z[7]));
  CDN_bmux8 g26(.sel0 (ctl[0]), .data0 (in_0[6]), .data1 (in_1[6]),
       .sel1 (ctl[1]), .data2 (in_2[6]), .data3 (in_3[6]), .sel2
       (ctl[2]), .data4 (in_4[6]), .data5 (in_5[6]), .data6 (in_6[6]),
       .data7 (in_7[6]), .z (z[6]));
  CDN_bmux8 g27(.sel0 (ctl[0]), .data0 (in_0[5]), .data1 (in_1[5]),
       .sel1 (ctl[1]), .data2 (in_2[5]), .data3 (in_3[5]), .sel2
       (ctl[2]), .data4 (in_4[5]), .data5 (in_5[5]), .data6 (in_6[5]),
       .data7 (in_7[5]), .z (z[5]));
  CDN_bmux8 g28(.sel0 (ctl[0]), .data0 (in_0[4]), .data1 (in_1[4]),
       .sel1 (ctl[1]), .data2 (in_2[4]), .data3 (in_3[4]), .sel2
       (ctl[2]), .data4 (in_4[4]), .data5 (in_5[4]), .data6 (in_6[4]),
       .data7 (in_7[4]), .z (z[4]));
  CDN_bmux8 g29(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .sel2
       (ctl[2]), .data4 (in_4[3]), .data5 (in_5[3]), .data6 (in_6[3]),
       .data7 (in_7[3]), .z (z[3]));
  CDN_bmux8 g30(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .sel2
       (ctl[2]), .data4 (in_4[2]), .data5 (in_5[2]), .data6 (in_6[2]),
       .data7 (in_7[2]), .z (z[2]));
  CDN_bmux8 g31(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .sel2
       (ctl[2]), .data4 (in_4[1]), .data5 (in_5[1]), .data6 (in_6[1]),
       .data7 (in_7[1]), .z (z[1]));
  CDN_bmux8 g32(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .sel2
       (ctl[2]), .data4 (in_4[0]), .data5 (in_5[0]), .data6 (in_6[0]),
       .data7 (in_7[0]), .z (z[0]));
endmodule

module fx68k_mux_2428(ctl, in_0, in_1, z);
  input [1:0] ctl;
  input [7:0] in_0, in_1;
  output [7:0] z;
  wire [1:0] ctl;
  wire [7:0] in_0, in_1;
  wire [7:0] z;
  CDN_mux2 g1(.sel0 (ctl[1]), .data0 (in_0[7]), .sel1 (ctl[0]), .data1
       (in_1[7]), .z (z[7]));
  CDN_mux2 g9(.sel0 (ctl[1]), .data0 (in_0[6]), .sel1 (ctl[0]), .data1
       (in_1[6]), .z (z[6]));
  CDN_mux2 g10(.sel0 (ctl[1]), .data0 (in_0[5]), .sel1 (ctl[0]), .data1
       (in_1[5]), .z (z[5]));
  CDN_mux2 g11(.sel0 (ctl[1]), .data0 (in_0[4]), .sel1 (ctl[0]), .data1
       (in_1[4]), .z (z[4]));
  CDN_mux2 g12(.sel0 (ctl[1]), .data0 (in_0[3]), .sel1 (ctl[0]), .data1
       (in_1[3]), .z (z[3]));
  CDN_mux2 g13(.sel0 (ctl[1]), .data0 (in_0[2]), .sel1 (ctl[0]), .data1
       (in_1[2]), .z (z[2]));
  CDN_mux2 g14(.sel0 (ctl[1]), .data0 (in_0[1]), .sel1 (ctl[0]), .data1
       (in_1[1]), .z (z[1]));
  CDN_mux2 g15(.sel0 (ctl[1]), .data0 (in_0[0]), .sel1 (ctl[0]), .data1
       (in_1[0]), .z (z[0]));
endmodule

module fx68k_excUnit(\Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] ,
     \Clks[extReset] , \Clks[clk] , enT1, enT2, enT3, enT4,
     \Nanod[abdIsByte] , \Nanod[dblDbh] , \Nanod[dblDbd] ,
     \Nanod[ablAbh] , \Nanod[ablAbd] , \Nanod[extAbh] , \Nanod[extDbh]
     , \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] , \Nanod[au2Pc] ,
     \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd] , \Nanod[alu2Dbd]
     , \Nanod[abd2Alub] , \Nanod[dbd2Alub] , \Nanod[alue2Dbd] ,
     \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] , \Nanod[abd2Dcr] ,
     \Nanod[aluFinish] , \Nanod[aluInit] , \Nanod[aluActrl] ,
     \Nanod[aluDctrl] , \Nanod[aluColumn] , \Nanod[rxlDbl] , \Nanod[rz]
     , \Nanod[abl2ryl] , \Nanod[dbl2ryl] , \Nanod[ryh2abh] ,
     \Nanod[ryh2dbh] , \Nanod[ryl2ab] , \Nanod[ryl2db] ,
     \Nanod[abh2ryh] , \Nanod[dbh2ryh] , \Nanod[abh2rxh] ,
     \Nanod[abl2rxl] , \Nanod[rxl2ab] , \Nanod[rxl2db] ,
     \Nanod[dbh2rxh] , \Nanod[dbl2rxl] , \Nanod[rxh2abh] ,
     \Nanod[rxh2dbh] , \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl]
     , \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
     , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
     \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
     \Nanod[dobCtrl] , \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob]
     , \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
     \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
     \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
     \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] , \Nanod[auCntrl]
     , \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
     \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
     \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
     \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
     \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
     \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
     \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
     \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
     \Nanod[waitBusFinish] , \Nanod[permStart] , \Irdecod[inhibitCcr] ,
     \Irdecod[macroTvn] , \Irdecod[ftuConst] , \Irdecod[ryIsAreg] ,
     \Irdecod[rxIsAreg] , \Irdecod[ry] , \Irdecod[rx] ,
     \Irdecod[isMovep] , \Irdecod[isByte] , \Irdecod[movemPreDecr] ,
     \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] ,
     \Irdecod[rxIsDt] , \Irdecod[toCcr] , \Irdecod[implicitSp] ,
     \Irdecod[isTas] , \Irdecod[isPcRel] , Ird, pswS, ftu, iEdb, ccr,
     alue, prenEmpty, au05z, dcr4, ze, aob0, AblOut, Irc, oEdb, eab);
  input \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset]
       , \Clks[clk] , enT1, enT2, enT3, enT4, \Nanod[abdIsByte] ,
       \Nanod[dblDbh] , \Nanod[dblDbd] , \Nanod[ablAbh] ,
       \Nanod[ablAbd] , \Nanod[extAbh] , \Nanod[extDbh] ,
       \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] , \Nanod[au2Pc] ,
       \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd] ,
       \Nanod[alu2Dbd] , \Nanod[abd2Alub] , \Nanod[dbd2Alub] ,
       \Nanod[alue2Dbd] , \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] ,
       \Nanod[abd2Dcr] , \Nanod[aluFinish] , \Nanod[aluInit] ,
       \Nanod[aluActrl] , \Nanod[rxlDbl] , \Nanod[rz] , \Nanod[abl2ryl]
       , \Nanod[dbl2ryl] , \Nanod[ryh2abh] , \Nanod[ryh2dbh] ,
       \Nanod[ryl2ab] , \Nanod[ryl2db] , \Nanod[abh2ryh] ,
       \Nanod[dbh2ryh] , \Nanod[abh2rxh] , \Nanod[abl2rxl] ,
       \Nanod[rxl2ab] , \Nanod[rxl2db] , \Nanod[dbh2rxh] ,
       \Nanod[dbl2rxl] , \Nanod[rxh2abh] , \Nanod[rxh2dbh] ,
       \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl] ,
       \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
       , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
       \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
       \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob] ,
       \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
       \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
       \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
       \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] ,
       \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
       \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
       \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
       \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
       \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
       \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
       \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
       \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
       \Nanod[waitBusFinish] , \Nanod[permStart] , \Irdecod[inhibitCcr]
       , \Irdecod[ryIsAreg] , \Irdecod[rxIsAreg] , \Irdecod[isMovep] ,
       \Irdecod[isByte] , \Irdecod[movemPreDecr] , \Irdecod[rxIsMovem]
       , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] , \Irdecod[rxIsDt] ,
       \Irdecod[toCcr] , \Irdecod[implicitSp] , \Irdecod[isTas] ,
       \Irdecod[isPcRel] , pswS;
  input [1:0] \Nanod[aluDctrl] , \Nanod[dobCtrl] ;
  input [2:0] \Nanod[aluColumn] , \Nanod[auCntrl] , \Irdecod[ry] ,
       \Irdecod[rx] ;
  input [5:0] \Irdecod[macroTvn] ;
  input [15:0] \Irdecod[ftuConst] , Ird, ftu, iEdb;
  output [7:0] ccr;
  output [15:0] alue, AblOut, Irc, oEdb;
  output prenEmpty, au05z, dcr4, ze, aob0;
  output [23:1] eab;
  wire \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset] ,
       \Clks[clk] , enT1, enT2, enT3, enT4, \Nanod[abdIsByte] ,
       \Nanod[dblDbh] , \Nanod[dblDbd] , \Nanod[ablAbh] ,
       \Nanod[ablAbd] , \Nanod[extAbh] , \Nanod[extDbh] ,
       \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] , \Nanod[au2Pc] ,
       \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd] ,
       \Nanod[alu2Dbd] , \Nanod[abd2Alub] , \Nanod[dbd2Alub] ,
       \Nanod[alue2Dbd] , \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] ,
       \Nanod[abd2Dcr] , \Nanod[aluFinish] , \Nanod[aluInit] ,
       \Nanod[aluActrl] , \Nanod[rxlDbl] , \Nanod[rz] , \Nanod[abl2ryl]
       , \Nanod[dbl2ryl] , \Nanod[ryh2abh] , \Nanod[ryh2dbh] ,
       \Nanod[ryl2ab] , \Nanod[ryl2db] , \Nanod[abh2ryh] ,
       \Nanod[dbh2ryh] , \Nanod[abh2rxh] , \Nanod[abl2rxl] ,
       \Nanod[rxl2ab] , \Nanod[rxl2db] , \Nanod[dbh2rxh] ,
       \Nanod[dbl2rxl] , \Nanod[rxh2abh] , \Nanod[rxh2dbh] ,
       \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl] ,
       \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
       , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
       \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
       \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob] ,
       \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
       \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
       \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
       \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] ,
       \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
       \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
       \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
       \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
       \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
       \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
       \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
       \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
       \Nanod[waitBusFinish] , \Nanod[permStart] , \Irdecod[inhibitCcr]
       , \Irdecod[ryIsAreg] , \Irdecod[rxIsAreg] , \Irdecod[isMovep] ,
       \Irdecod[isByte] , \Irdecod[movemPreDecr] , \Irdecod[rxIsMovem]
       , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] , \Irdecod[rxIsDt] ,
       \Irdecod[toCcr] , \Irdecod[implicitSp] , \Irdecod[isTas] ,
       \Irdecod[isPcRel] , pswS;
  wire [1:0] \Nanod[aluDctrl] , \Nanod[dobCtrl] ;
  wire [2:0] \Nanod[aluColumn] , \Nanod[auCntrl] , \Irdecod[ry] ,
       \Irdecod[rx] ;
  wire [5:0] \Irdecod[macroTvn] ;
  wire [15:0] \Irdecod[ftuConst] , Ird, ftu, iEdb;
  wire [7:0] ccr;
  wire [15:0] alue, AblOut, Irc, oEdb;
  wire prenEmpty, au05z, dcr4, ze, aob0;
  wire [23:1] eab;
  wire [15:0] prenLatch;
  wire [3:0] prHbit;
  wire [3:0] dcrInput;
  wire [15:0] dcrCode;
  wire [15:0] dobInput;
  wire [15:0] dbin;
  wire [15:0] alub;
  wire [15:0] Dbd;
  wire [15:0] Abd;
  wire [15:0] aluOut;
  wire [3:0] rxReg;
  wire [3:0] ryReg;
  wire [4:0] rxMux;
  wire [4:0] ryMux;
  wire [15:0] Dbh;
  wire [15:0] Dbl;
  wire [31:0] auInpMux;
  wire [3:0] movemRx;
  wire [31:0] auReg;
  wire [4:0] actualRx;
  wire [15:0] \regs68L[0] ;
  wire [15:0] \regs68L[1] ;
  wire [15:0] \regs68L[2] ;
  wire [15:0] \regs68L[3] ;
  wire [15:0] \regs68L[4] ;
  wire [15:0] \regs68L[5] ;
  wire [15:0] \regs68L[6] ;
  wire [15:0] \regs68L[7] ;
  wire [15:0] \regs68L[8] ;
  wire [15:0] \regs68L[9] ;
  wire [15:0] \regs68L[10] ;
  wire [15:0] \regs68L[11] ;
  wire [15:0] \regs68L[12] ;
  wire [15:0] \regs68L[13] ;
  wire [15:0] \regs68L[14] ;
  wire [15:0] \regs68L[15] ;
  wire [15:0] \regs68L[16] ;
  wire [15:0] \regs68L[17] ;
  wire [4:0] actualRy;
  wire [15:0] PcL;
  wire [15:0] Atl;
  wire [15:0] ablMux;
  wire [15:0] \regs68L[actualRy] ;
  wire [15:0] \regs68L[actualRx] ;
  wire [15:0] Abh;
  wire [15:0] \regs68H[0] ;
  wire [15:0] \regs68H[1] ;
  wire [15:0] \regs68H[2] ;
  wire [15:0] \regs68H[3] ;
  wire [15:0] \regs68H[4] ;
  wire [15:0] \regs68H[5] ;
  wire [15:0] \regs68H[6] ;
  wire [15:0] \regs68H[7] ;
  wire [15:0] \regs68H[8] ;
  wire [15:0] \regs68H[9] ;
  wire [15:0] \regs68H[10] ;
  wire [15:0] \regs68H[11] ;
  wire [15:0] \regs68H[12] ;
  wire [15:0] \regs68H[13] ;
  wire [15:0] \regs68H[14] ;
  wire [15:0] \regs68H[15] ;
  wire [15:0] \regs68H[16] ;
  wire [15:0] \regs68H[17] ;
  wire [15:0] \regs68H[actualRx] ;
  wire [15:0] \regs68H[actualRy] ;
  wire [15:0] Ath;
  wire [15:0] PcH;
  wire [15:0] dbhMux;
  wire [31:0] aob;
  wire [15:0] abhMux;
  wire [15:0] abdMux;
  wire [15:0] preAbl;
  wire [15:0] preAbh;
  wire [15:0] preAbd;
  wire [15:0] dblMux;
  wire [15:0] preDbd;
  wire [15:0] preDbh;
  wire [15:0] preDbl;
  wire [15:0] dcrOutput;
  wire [15:0] dbdMux;
  wire [15:0] Abl;
  wire Pch2Abh, Pch2Dbh, Pcl2Abl, Pcl2Dbl, UNCONNECTED442,
       UNCONNECTED443, UNCONNECTED444, UNCONNECTED445;
  wire UNCONNECTED446, UNCONNECTED447, UNCONNECTED448, UNCONNECTED449,
       UNCONNECTED450, UNCONNECTED451, UNCONNECTED452, UNCONNECTED453;
  wire UNCONNECTED454, UNCONNECTED455, UNCONNECTED456, UNCONNECTED457,
       UNCONNECTED458, UNCONNECTED459, UNCONNECTED460, UNCONNECTED461;
  wire UNCONNECTED462, UNCONNECTED463, UNCONNECTED464, UNCONNECTED465,
       UNCONNECTED466, UNCONNECTED467, UNCONNECTED468, UNCONNECTED469;
  wire UNCONNECTED470, UNCONNECTED471, UNCONNECTED472, UNCONNECTED473,
       UNCONNECTED474, UNCONNECTED475, UNCONNECTED476, UNCONNECTED477;
  wire UNCONNECTED478, UNCONNECTED479, UNCONNECTED480, UNCONNECTED481,
       UNCONNECTED482, _X_, abdIdle, abdIsByte;
  wire abh2Pch, abhIdle, abl2Pcl, ablIdle, alueClkEn, au2Aob,
       byteNotSpAlign, dbdIdle;
  wire dbh2Pch, dbhIdle, dbl2Pcl, dblIdle, dobIdle, n_6, n_8, n_9;
  wire n_10, n_11, n_13, n_15, n_16, n_17, n_18, n_19;
  wire n_20, n_28, n_29, n_30, n_32, n_33, n_34, n_36;
  wire n_37, n_38, n_62, n_76, n_90, n_118, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_423, n_424, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_449, n_451, n_453, n_456;
  wire n_457, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_483, n_484, n_485;
  wire n_486, n_492, n_493, n_494, n_495, n_501, n_502, n_503;
  wire n_505, n_517, n_518, n_520, n_521, n_523, n_524, n_525;
  wire n_535, n_536, n_537, n_551, n_552, n_553, n_554, n_555;
  wire n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_590, n_591, n_593, n_594, n_596, n_597, n_599, n_600;
  wire n_602, n_603, n_605, n_606, n_608, n_609, n_611, n_612;
  wire n_614, n_615, n_617, n_618, n_620, n_621, n_623, n_624;
  wire n_626, n_627, n_629, n_630, n_632, n_633, n_635, n_636;
  wire n_639, n_641, n_643, n_644, n_653, n_654, n_666, n_667;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
  wire n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708;
  wire n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716;
  wire n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724;
  wire n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732;
  wire n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740;
  wire n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756;
  wire n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764;
  wire n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780;
  wire n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788;
  wire n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796;
  wire n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804;
  wire n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820;
  wire n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900;
  wire n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964;
  wire n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972;
  wire n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980;
  wire n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988;
  wire n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996;
  wire n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004;
  wire n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012;
  wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1027, n_1028, n_1029, n_1030;
  wire n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038;
  wire n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046;
  wire n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054;
  wire n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062;
  wire n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070;
  wire n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078;
  wire n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086;
  wire n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094;
  wire n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102;
  wire n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134;
  wire n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1153, n_1154, n_1155, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186;
  wire n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194;
  wire n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202;
  wire n_1203, n_1204, n_1205, n_1206, n_1207, n_1209, n_1210, n_1211;
  wire n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219;
  wire n_1220, n_1221, n_1222, n_1223, n_1224, n_1226, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264;
  wire n_1265, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292;
  wire n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300;
  wire n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308;
  wire n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316;
  wire n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1344, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362;
  wire n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370;
  wire n_1371, n_1372, n_1373, n_1374, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387;
  wire n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395;
  wire n_1396, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413;
  wire n_1414, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425;
  wire n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433;
  wire n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441;
  wire n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465;
  wire n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473;
  wire n_1474, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483;
  wire n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491;
  wire n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499;
  wire n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523;
  wire n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531;
  wire n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539;
  wire n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547;
  wire n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555;
  wire n_1556, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565;
  wire n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573;
  wire n_1574, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585;
  wire n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593;
  wire n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601;
  wire n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609;
  wire n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617;
  wire n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625;
  wire n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633;
  wire n_1634, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643;
  wire n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651;
  wire n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683;
  wire n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691;
  wire n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699;
  wire n_1700, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729;
  wire n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737;
  wire n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745;
  wire n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753;
  wire n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761;
  wire n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769;
  wire n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777;
  wire n_1778, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787;
  wire n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795;
  wire n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803;
  wire n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811;
  wire n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819;
  wire n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827;
  wire n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835;
  wire n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843;
  wire n_1844, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853;
  wire n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861;
  wire n_1862, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873;
  wire n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881;
  wire n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889;
  wire n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897;
  wire n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905;
  wire n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913;
  wire n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921;
  wire n_1922, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931;
  wire n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939;
  wire n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947;
  wire n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955;
  wire n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963;
  wire n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971;
  wire n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979;
  wire n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987;
  wire n_1988, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997;
  wire n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005;
  wire n_2006, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017;
  wire n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025;
  wire n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033;
  wire n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057;
  wire n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065;
  wire n_2066, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075;
  wire n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083;
  wire n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091;
  wire n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099;
  wire n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107;
  wire n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115;
  wire n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123;
  wire n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131;
  wire n_2132, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141;
  wire n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149;
  wire n_2150, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161;
  wire n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169;
  wire n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177;
  wire n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185;
  wire n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193;
  wire n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201;
  wire n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209;
  wire n_2210, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219;
  wire n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227;
  wire n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235;
  wire n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243;
  wire n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251;
  wire n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259;
  wire n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267;
  wire n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275;
  wire n_2276, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285;
  wire n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293;
  wire n_2294, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305;
  wire n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313;
  wire n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321;
  wire n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329;
  wire n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337;
  wire n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345;
  wire n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353;
  wire n_2354, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363;
  wire n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371;
  wire n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379;
  wire n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387;
  wire n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395;
  wire n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403;
  wire n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411;
  wire n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419;
  wire n_2420, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429;
  wire n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437;
  wire n_2438, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449;
  wire n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457;
  wire n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465;
  wire n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473;
  wire n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481;
  wire n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489;
  wire n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497;
  wire n_2498, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507;
  wire n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515;
  wire n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523;
  wire n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531;
  wire n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539;
  wire n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547;
  wire n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555;
  wire n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563;
  wire n_2564, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573;
  wire n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581;
  wire n_2582, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593;
  wire n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601;
  wire n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609;
  wire n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617;
  wire n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625;
  wire n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633;
  wire n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641;
  wire n_2642, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651;
  wire n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659;
  wire n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667;
  wire n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675;
  wire n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683;
  wire n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
  wire n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699;
  wire n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707;
  wire n_2708, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717;
  wire n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725;
  wire n_2726, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737;
  wire n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745;
  wire n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753;
  wire n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761;
  wire n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769;
  wire n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777;
  wire n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785;
  wire n_2786, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795;
  wire n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803;
  wire n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811;
  wire n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819;
  wire n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827;
  wire n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835;
  wire n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843;
  wire n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851;
  wire n_2852, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861;
  wire n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869;
  wire n_2870, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881;
  wire n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889;
  wire n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905;
  wire n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913;
  wire n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921;
  wire n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929;
  wire n_2930, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939;
  wire n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947;
  wire n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955;
  wire n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963;
  wire n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971;
  wire n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979;
  wire n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987;
  wire n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995;
  wire n_2996, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005;
  wire n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013;
  wire n_3014, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025;
  wire n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033;
  wire n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041;
  wire n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049;
  wire n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057;
  wire n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065;
  wire n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073;
  wire n_3074, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083;
  wire n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091;
  wire n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099;
  wire n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107;
  wire n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115;
  wire n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123;
  wire n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131;
  wire n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139;
  wire n_3140, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149;
  wire n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157;
  wire n_3158, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169;
  wire n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177;
  wire n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185;
  wire n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193;
  wire n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201;
  wire n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209;
  wire n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217;
  wire n_3218, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227;
  wire n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235;
  wire n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243;
  wire n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251;
  wire n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259;
  wire n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267;
  wire n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275;
  wire n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283;
  wire n_3284, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293;
  wire n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301;
  wire n_3302, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313;
  wire n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321;
  wire n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329;
  wire n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337;
  wire n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345;
  wire n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353;
  wire n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361;
  wire n_3362, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371;
  wire n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379;
  wire n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387;
  wire n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395;
  wire n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403;
  wire n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411;
  wire n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419;
  wire n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427;
  wire n_3428, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437;
  wire n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445;
  wire n_3446, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457;
  wire n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465;
  wire n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473;
  wire n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481;
  wire n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489;
  wire n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497;
  wire n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505;
  wire n_3506, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515;
  wire n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523;
  wire n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531;
  wire n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539;
  wire n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547;
  wire n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555;
  wire n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563;
  wire n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571;
  wire n_3572, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581;
  wire n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589;
  wire n_3590, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601;
  wire n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609;
  wire n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617;
  wire n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625;
  wire n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633;
  wire n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641;
  wire n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649;
  wire n_3650, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659;
  wire n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667;
  wire n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675;
  wire n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683;
  wire n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691;
  wire n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699;
  wire n_3700, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723;
  wire n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731;
  wire n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739;
  wire n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747;
  wire n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755;
  wire n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763;
  wire n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771;
  wire n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779;
  wire n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787;
  wire n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795;
  wire n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803;
  wire n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811;
  wire n_3812, n_3813, n_3814, n_3817, n_3818, n_3819, n_3820, n_3821;
  wire n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829;
  wire n_3830, n_3831, n_3832, n_3837, n_3838, n_3839, n_3840, n_3841;
  wire n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849;
  wire n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857;
  wire n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865;
  wire n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873;
  wire n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881;
  wire n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889;
  wire n_3890, n_3891, n_3892, n_3895, n_3896, n_3897, n_3898, n_3899;
  wire n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907;
  wire n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915;
  wire n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923;
  wire n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, n_3931;
  wire n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939;
  wire n_3940, n_3941, n_3942, n_3945, n_3946, n_3947, n_3948, n_3949;
  wire n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957;
  wire n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965;
  wire n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973;
  wire n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981;
  wire n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989;
  wire n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997;
  wire n_3998, n_3999, n_4000, n_4003, n_4004, n_4005, n_4006, n_4007;
  wire n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015;
  wire n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023;
  wire n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031;
  wire n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039;
  wire n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047;
  wire n_4048, n_4049, n_4050, n_4178, n_4179, n_4181, n_4182, n_4183;
  wire n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191;
  wire n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199;
  wire n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207;
  wire n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215;
  wire n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223;
  wire n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231;
  wire n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239;
  wire n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247;
  wire n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255;
  wire n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263;
  wire n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271;
  wire n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279;
  wire n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287;
  wire n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295;
  wire n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303;
  wire n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311;
  wire n_4312, n_4313, n_4314, n_4315, n_4318, n_4319, n_4320, n_4321;
  wire n_4322, n_4323, n_4324, n_4326, n_4327, n_4328, n_4331, n_4332;
  wire n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341;
  wire n_4342, n_4350, n_4351, n_4353, n_4354, n_4355, n_4356, n_4357;
  wire n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4368, n_4369;
  wire n_4371, n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378;
  wire n_4379, n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386;
  wire n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394;
  wire n_4395, n_4396, n_4397, n_4398, n_4399, n_4400, n_4403, n_4404;
  wire n_4405, n_4406, n_4407, n_4409, n_4410, n_4411, n_4413, n_4414;
  wire n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423;
  wire n_4424, n_4432, n_4433, n_4435, n_4436, n_4437, n_4438, n_4439;
  wire n_4440, n_4441, n_4442, n_4443, n_4444, n_4448, n_4449, n_4451;
  wire n_4452, n_4453, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459;
  wire n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467;
  wire n_4468, n_4469, n_4470, n_4471, n_4472, n_4473, n_4474, n_4475;
  wire n_4476, n_4477, n_4478, n_4479, n_4482, n_4483, n_4484, n_4485;
  wire n_4486, n_4488, n_4489, n_4490, n_4492, n_4493, n_4495, n_4496;
  wire n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4511;
  wire n_4512, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520;
  wire n_4521, n_4522, n_4523, n_4527, n_4528, n_4530, n_4531, n_4532;
  wire n_4533, n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540;
  wire n_4541, n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548;
  wire n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556;
  wire n_4557, n_4558, n_4561, n_4562, n_4563, n_4564, n_4565, n_4567;
  wire n_4568, n_4569, n_4571, n_4572, n_4574, n_4575, n_4576, n_4577;
  wire n_4578, n_4579, n_4580, n_4581, n_4582, n_4590, n_4591, n_4593;
  wire n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601;
  wire n_4602, n_4606, n_4607, n_4609, n_4610, n_4611, n_4612, n_4613;
  wire n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621;
  wire n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629;
  wire n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637;
  wire n_4640, n_4641, n_4642, n_4643, n_4644, n_4646, n_4647, n_4648;
  wire n_4650, n_4651, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658;
  wire n_4659, n_4660, n_4661, n_4669, n_4670, n_4672, n_4673, n_4674;
  wire n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4685;
  wire n_4686, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693, n_4694;
  wire n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701, n_4702;
  wire n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709, n_4710;
  wire n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4719, n_4720;
  wire n_4721, n_4722, n_4723, n_4725, n_4726, n_4727, n_4729, n_4730;
  wire n_4732, n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739;
  wire n_4740, n_4748, n_4749, n_4751, n_4752, n_4753, n_4754, n_4755;
  wire n_4756, n_4757, n_4758, n_4759, n_4760, n_4764, n_4765, n_4767;
  wire n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775;
  wire n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783;
  wire n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791;
  wire n_4792, n_4793, n_4794, n_4795, n_4798, n_4799, n_4800, n_4801;
  wire n_4802, n_4804, n_4805, n_4806, n_4808, n_4809, n_4811, n_4812;
  wire n_4813, n_4814, n_4815, n_4816, n_4817, n_4818, n_4819, n_4827;
  wire n_4828, n_4830, n_4831, n_4832, n_4833, n_4834, n_4835, n_4836;
  wire n_4837, n_4838, n_4839, n_4843, n_4844, n_4846, n_4847, n_4848;
  wire n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856;
  wire n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864;
  wire n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872;
  wire n_4873, n_4874, n_4877, n_4878, n_4879, n_4880, n_4881, n_4883;
  wire n_4884, n_4885, n_4887, n_4888, n_4890, n_4891, n_4892, n_4893;
  wire n_4894, n_4895, n_4896, n_4897, n_4898, n_4906, n_4907, n_4909;
  wire n_4910, n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917;
  wire n_4918, n_4922, n_4923, n_4925, n_4926, n_4927, n_4928, n_4929;
  wire n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937;
  wire n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945;
  wire n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953;
  wire n_4956, n_4957, n_4958, n_4959, n_4960, n_4962, n_4963, n_4964;
  wire n_4966, n_4967, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974;
  wire n_4975, n_4976, n_4977, n_4985, n_4986, n_4988, n_4989, n_4990;
  wire n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_5001;
  wire n_5002, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010;
  wire n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018;
  wire n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026;
  wire n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, n_5035, n_5036;
  wire n_5037, n_5038, n_5039, n_5041, n_5042, n_5043, n_5045, n_5046;
  wire n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055;
  wire n_5056, n_5064, n_5065, n_5067, n_5068, n_5069, n_5070, n_5071;
  wire n_5072, n_5073, n_5074, n_5075, n_5076, n_5080, n_5081, n_5083;
  wire n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091;
  wire n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099;
  wire n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107;
  wire n_5108, n_5109, n_5110, n_5111, n_5114, n_5115, n_5116, n_5117;
  wire n_5118, n_5120, n_5121, n_5122, n_5124, n_5125, n_5127, n_5128;
  wire n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5143;
  wire n_5144, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152;
  wire n_5153, n_5154, n_5155, n_5159, n_5160, n_5162, n_5163, n_5164;
  wire n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172;
  wire n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180;
  wire n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5188;
  wire n_5189, n_5190, n_5193, n_5194, n_5195, n_5196, n_5197, n_5199;
  wire n_5200, n_5201, n_5203, n_5204, n_5206, n_5207, n_5208, n_5209;
  wire n_5210, n_5211, n_5212, n_5213, n_5214, n_5222, n_5223, n_5225;
  wire n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232, n_5233;
  wire n_5234, n_5238, n_5239, n_5241, n_5242, n_5243, n_5244, n_5245;
  wire n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252, n_5253;
  wire n_5254, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260, n_5261;
  wire n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269;
  wire n_5272, n_5273, n_5274, n_5275, n_5276, n_5278, n_5279, n_5280;
  wire n_5282, n_5283, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290;
  wire n_5291, n_5292, n_5293, n_5301, n_5302, n_5304, n_5305, n_5306;
  wire n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313, n_5317;
  wire n_5318, n_5320, n_5321, n_5322, n_5323, n_5324, n_5325, n_5326;
  wire n_5327, n_5328, n_5329, n_5330, n_5331, n_5332, n_5333, n_5334;
  wire n_5335, n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342;
  wire n_5343, n_5344, n_5345, n_5346, n_5347, n_5348, n_5351, n_5352;
  wire n_5353, n_5354, n_5355, n_5357, n_5358, n_5359, n_5361, n_5362;
  wire n_5364, n_5365, n_5366, n_5367, n_5368, n_5369, n_5370, n_5371;
  wire n_5372, n_5380, n_5381, n_5383, n_5384, n_5385, n_5386, n_5387;
  wire n_5388, n_5389, n_5390, n_5391, n_5392, n_5396, n_5397, n_5399;
  wire n_5400, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407;
  wire n_5408, n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415;
  wire n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423;
  wire n_5424, n_5425, n_5426, n_5427, n_5430, n_5431, n_5432, n_5433;
  wire n_5434, n_5436, n_5437, n_5438, n_5440, n_5441, n_5443, n_5444;
  wire n_5445, n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5459;
  wire n_5460, n_5462, n_5463, n_5464, n_5465, n_5466, n_5467, n_5468;
  wire n_5469, n_5470, n_5471, n_5475, n_5476, n_5478, n_5479, n_5480;
  wire n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488;
  wire n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496;
  wire n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504;
  wire n_5505, n_5506, n_5509, n_5510, n_5511, n_5512, n_5513, n_5515;
  wire n_5516, n_5517, n_5519, n_5520, n_5522, n_5523, n_5524, n_5525;
  wire n_5526, n_5527, n_5528, n_5529, n_5530, n_5538, n_5539, n_5541;
  wire n_5542, n_5543, n_5544, n_5545, n_5546, n_5547, n_5548, n_5549;
  wire n_5550, n_5554, n_5555, n_5557, n_5558, n_5559, n_5560, n_5561;
  wire n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, n_5569;
  wire n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576, n_5577;
  wire n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585;
  wire n_5588, n_5589, n_5590, n_5591, n_5592, n_5594, n_5595, n_5596;
  wire n_5598, n_5599, n_5601, n_5602, n_5603, n_5604, n_5605, n_5606;
  wire n_5607, n_5608, n_5609, n_5617, n_5618, n_5620, n_5621, n_5622;
  wire n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629, n_5633;
  wire n_5634, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641, n_5642;
  wire n_5643, n_5644, n_5645, n_5646, n_5647, n_5648, n_5649, n_5650;
  wire n_5651, n_5652, n_5653, n_5654, n_5655, n_5656, n_5657, n_5658;
  wire n_5659, n_5660, n_5661, n_5662, n_5663, n_5664, n_5667, n_5668;
  wire n_5669, n_5670, n_5671, n_5673, n_5674, n_5675, n_5677, n_5678;
  wire n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686, n_5687;
  wire n_5688, n_5696, n_5697, n_5699, n_5700, n_5701, n_5702, n_5703;
  wire n_5704, n_5705, n_5706, n_5707, n_5708, n_5712, n_5713, n_5715;
  wire n_5716, n_5717, n_5718, n_5719, n_5720, n_5721, n_5722, n_5723;
  wire n_5724, n_5725, n_5726, n_5727, n_5728, n_5729, n_5730, n_5731;
  wire n_5732, n_5733, n_5734, n_5735, n_5736, n_5737, n_5738, n_5739;
  wire n_5740, n_5741, n_5742, n_5744, n_5745, n_5746, n_5747, n_5748;
  wire n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5756;
  wire n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764;
  wire n_5765, n_5766, n_5767, n_5769, n_5770, n_5771, n_5772, n_5773;
  wire n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780, n_5781;
  wire n_5782, n_5783, n_5784, n_5785, n_5786, n_5787, n_5788, n_5789;
  wire n_5790, n_5791, n_5793, n_5794, n_5795, n_5796, n_5797, n_5798;
  wire n_5799, n_5800, n_5801, n_5802, n_5803, n_5804, n_5805, n_5806;
  wire n_5807, n_5808, n_5809, n_5810, n_5811, n_5812, n_5813, n_5814;
  wire n_5815, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822, n_5823;
  wire n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831;
  wire n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838, n_5839;
  wire n_5841, n_5842, n_5843, n_5844, n_5845, n_5846, n_5847, n_5848;
  wire n_5849, n_5850, n_5851, n_5852, n_5853, n_5854, n_5855, n_5856;
  wire n_5857, n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5865;
  wire n_5866, n_5867, n_5868, n_5869, n_5870, n_5871, n_5872, n_5873;
  wire n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880, n_5881;
  wire n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5889, n_5890;
  wire n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898;
  wire n_5899, n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906;
  wire n_5907, n_5908, n_5909, n_5910, n_5911, n_5913, n_5914, n_5915;
  wire n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923;
  wire n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931;
  wire n_5932, n_5933, n_5934, n_5935, n_5937, n_5938, n_5939, n_5940;
  wire n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948;
  wire n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956;
  wire n_5957, n_5958, n_5959, n_5961, n_5962, n_5963, n_5964, n_5965;
  wire n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972, n_5973;
  wire n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980, n_5981;
  wire n_5982, n_5983, n_5985, n_5986, n_5987, n_5988, n_5989, n_5990;
  wire n_5991, n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998;
  wire n_5999, n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6006;
  wire n_6007, n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015;
  wire n_6016, n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023;
  wire n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031;
  wire n_6033, n_6034, n_6035, n_6036, n_6037, n_6038, n_6039, n_6040;
  wire n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048;
  wire n_6049, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6057;
  wire n_6058, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064, n_6065;
  wire n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072, n_6073;
  wire n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6081, n_6082;
  wire n_6083, n_6084, n_6085, n_6086, n_6087, n_6088, n_6089, n_6090;
  wire n_6091, n_6092, n_6093, n_6094, n_6095, n_6096, n_6097, n_6098;
  wire n_6099, n_6100, n_6101, n_6102, n_6103, n_6105, n_6106, n_6107;
  wire n_6108, n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, n_6115;
  wire n_6116, n_6117, n_6118, n_6119, n_6120, n_6121, n_6122, n_6123;
  wire n_6124, n_6125, n_6126, n_6127, n_6129, n_6130, n_6131, n_6132;
  wire n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139, n_6140;
  wire n_6141, n_6142, n_6143, n_6144, n_6145, n_6146, n_6147, n_6148;
  wire n_6149, n_6150, n_6151, n_6153, n_6154, n_6155, n_6156, n_6157;
  wire n_6158, n_6159, n_6160, n_6161, n_6162, n_6163, n_6164, n_6165;
  wire n_6166, n_6167, n_6168, n_6169, n_6170, n_6171, n_6172, n_6173;
  wire n_6174, n_6175, n_6176, n_6177, n_6178, n_6179, n_6180, n_6181;
  wire n_6182, n_6183, n_6184, n_6185, n_6186, n_6187, n_6188, n_6189;
  wire n_6190, n_6191, n_6192, n_6193, n_6194, n_6195, n_6196, n_6197;
  wire n_6198, n_6199, n_6200, n_6201, n_6202, n_6204, n_6205, n_6206;
  wire n_6207, n_6208, n_6209, n_6210, n_6211, n_6212, n_6213, n_6214;
  wire n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6222;
  wire n_6223, n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230;
  wire n_6231, n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238;
  wire n_6239, n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246;
  wire n_6247, n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254;
  wire n_6255, n_6256, n_6257, n_6258, n_6259, n_6260, n_6261, n_6262;
  wire n_6263, n_6264, n_6265, n_6266, n_6267, n_6269, n_6270, n_6271;
  wire n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279;
  wire n_6280, n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287;
  wire n_6288, n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295;
  wire n_6296, n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303;
  wire n_6304, n_6305, n_6306, n_6307, n_6349, n_6350, n_6351, n_6352;
  wire n_8229, n_8230, n_8231, n_8232, n_8233, n_8234, n_8235, n_8236;
  wire n_8237, n_8238, n_8239, n_8240, n_8241, n_8242, n_8243, n_8244;
  wire n_8245, n_8374, n_8375, n_8376, n_8377, n_8378, n_8379, n_8380;
  wire n_8381, n_8382, n_8384, n_8385, n_8386, n_8387, n_8388, n_8389;
  wire n_8390, n_8391, n_8392, n_8443, n_8444, n_8445, n_8502, n_8503;
  wire n_8504, n_8505, n_8506, n_8507, n_8616, n_8617, n_8618, rxIsAreg;
  wire rxIsSp, rxl2Abd, rxl2Abl, rxl2Dbd, rxl2Dbl, ryIsAreg, ryIsSp,
       ryl2Abd;
  wire ryl2Abl, ryl2Dbd, ryl2Dbl;
  fx68k_pren rmPren(.mask (prenLatch), .hbit (prHbit));
  fx68k_onehotEncoder4 dcrDecoder(.bin (dcrInput), .bitMap (dcrCode));
  fx68k_dataIo dataIo(.\Clks[enPhi2]  (\Clks[enPhi2] ), .\Clks[enPhi1] 
       (\Clks[enPhi1] ), .\Clks[pwrUp]  (\Clks[pwrUp] ),
       .\Clks[extReset]  (\Clks[extReset] ), .\Clks[clk]  (\Clks[clk]
       ), .enT1 (enT1), .enT2 (enT2), .enT3 (enT3), .enT4 (enT4),
       .\Nanod[abdIsByte]  (\Nanod[abdIsByte] ), .\Nanod[dblDbh] 
       (\Nanod[dblDbh] ), .\Nanod[dblDbd]  (\Nanod[dblDbd] ),
       .\Nanod[ablAbh]  (\Nanod[ablAbh] ), .\Nanod[ablAbd] 
       (\Nanod[ablAbd] ), .\Nanod[extAbh]  (\Nanod[extAbh] ),
       .\Nanod[extDbh]  (\Nanod[extDbh] ), .\Nanod[dbin2Dbd] 
       (\Nanod[dbin2Dbd] ), .\Nanod[dbin2Abd]  (\Nanod[dbin2Abd] ),
       .\Nanod[au2Pc]  (\Nanod[au2Pc] ), .\Nanod[au2Ab]  (\Nanod[au2Ab]
       ), .\Nanod[au2Db]  (\Nanod[au2Db] ), .\Nanod[alu2Abd] 
       (\Nanod[alu2Abd] ), .\Nanod[alu2Dbd]  (\Nanod[alu2Dbd] ),
       .\Nanod[abd2Alub]  (\Nanod[abd2Alub] ), .\Nanod[dbd2Alub] 
       (\Nanod[dbd2Alub] ), .\Nanod[alue2Dbd]  (\Nanod[alue2Dbd] ),
       .\Nanod[dbd2Alue]  (\Nanod[dbd2Alue] ), .\Nanod[dcr2Dbd] 
       (\Nanod[dcr2Dbd] ), .\Nanod[abd2Dcr]  (\Nanod[abd2Dcr] ),
       .\Nanod[aluFinish]  (\Nanod[aluFinish] ), .\Nanod[aluInit] 
       (\Nanod[aluInit] ), .\Nanod[aluActrl]  (\Nanod[aluActrl] ),
       .\Nanod[aluDctrl]  (\Nanod[aluDctrl] ), .\Nanod[aluColumn] 
       (\Nanod[aluColumn] ), .\Nanod[rxlDbl]  (\Nanod[rxlDbl] ),
       .\Nanod[rz]  (\Nanod[rz] ), .\Nanod[abl2ryl]  (\Nanod[abl2ryl]
       ), .\Nanod[dbl2ryl]  (\Nanod[dbl2ryl] ), .\Nanod[ryh2abh] 
       (\Nanod[ryh2abh] ), .\Nanod[ryh2dbh]  (\Nanod[ryh2dbh] ),
       .\Nanod[ryl2ab]  (\Nanod[ryl2ab] ), .\Nanod[ryl2db] 
       (\Nanod[ryl2db] ), .\Nanod[abh2ryh]  (\Nanod[abh2ryh] ),
       .\Nanod[dbh2ryh]  (\Nanod[dbh2ryh] ), .\Nanod[abh2rxh] 
       (\Nanod[abh2rxh] ), .\Nanod[abl2rxl]  (\Nanod[abl2rxl] ),
       .\Nanod[rxl2ab]  (\Nanod[rxl2ab] ), .\Nanod[rxl2db] 
       (\Nanod[rxl2db] ), .\Nanod[dbh2rxh]  (\Nanod[dbh2rxh] ),
       .\Nanod[dbl2rxl]  (\Nanod[dbl2rxl] ), .\Nanod[rxh2abh] 
       (\Nanod[rxh2abh] ), .\Nanod[rxh2dbh]  (\Nanod[rxh2dbh] ),
       .\Nanod[pchabh]  (\Nanod[pchabh] ), .\Nanod[pclabl] 
       (\Nanod[pclabl] ), .\Nanod[pcldbl]  (\Nanod[pcldbl] ),
       .\Nanod[pchdbh]  (\Nanod[pchdbh] ), .\Nanod[ssp]  (\Nanod[ssp]
       ), .\Nanod[reg2dbh]  (\Nanod[reg2dbh] ), .\Nanod[reg2dbl] 
       (\Nanod[reg2dbl] ), .\Nanod[dbl2reg]  (\Nanod[dbl2reg] ),
       .\Nanod[dbh2reg]  (\Nanod[dbh2reg] ), .\Nanod[reg2abh] 
       (\Nanod[reg2abh] ), .\Nanod[reg2abl]  (\Nanod[reg2abl] ),
       .\Nanod[abl2reg]  (\Nanod[abl2reg] ), .\Nanod[abh2reg] 
       (\Nanod[abh2reg] ), .\Nanod[dobCtrl]  (\Nanod[dobCtrl] ),
       .\Nanod[updSsw]  (\Nanod[updSsw] ), .\Nanod[aob2Ab] 
       (\Nanod[aob2Ab] ), .\Nanod[au2Aob]  (\Nanod[au2Aob] ),
       .\Nanod[ab2Aob]  (\Nanod[ab2Aob] ), .\Nanod[db2Aob] 
       (\Nanod[db2Aob] ), .\Nanod[ath2Abh]  (\Nanod[ath2Abh] ),
       .\Nanod[ath2Dbh]  (\Nanod[ath2Dbh] ), .\Nanod[dbh2Ath] 
       (\Nanod[dbh2Ath] ), .\Nanod[abh2Ath]  (\Nanod[abh2Ath] ),
       .\Nanod[atl2Dbl]  (\Nanod[atl2Dbl] ), .\Nanod[atl2Abl] 
       (\Nanod[atl2Abl] ), .\Nanod[abl2Atl]  (\Nanod[abl2Atl] ),
       .\Nanod[dbl2Atl]  (\Nanod[dbl2Atl] ), .\Nanod[toIrc] 
       (\Nanod[toIrc] ), .\Nanod[todbin]  (\Nanod[todbin] ),
       .\Nanod[auCntrl]  (\Nanod[auCntrl] ), .\Nanod[noSpAlign] 
       (\Nanod[noSpAlign] ), .\Nanod[auClkEn]  (\Nanod[auClkEn] ),
       .\Nanod[Ir2Ird]  (\Nanod[Ir2Ird] ), .\Nanod[initST] 
       (\Nanod[initST] ), .\Nanod[ssw2Ftu]  (\Nanod[ssw2Ftu] ),
       .\Nanod[ird2Ftu]  (\Nanod[ird2Ftu] ), .\Nanod[pswIToFtu] 
       (\Nanod[pswIToFtu] ), .\Nanod[ftu2Ccr]  (\Nanod[ftu2Ccr] ),
       .\Nanod[sr2Ftu]  (\Nanod[sr2Ftu] ), .\Nanod[ftu2Sr] 
       (\Nanod[ftu2Sr] ), .\Nanod[inl2psw]  (\Nanod[inl2psw] ),
       .\Nanod[updPren]  (\Nanod[updPren] ), .\Nanod[abl2Pren] 
       (\Nanod[abl2Pren] ), .\Nanod[ftu2Abl]  (\Nanod[ftu2Abl] ),
       .\Nanod[ftu2Dbl]  (\Nanod[ftu2Dbl] ), .\Nanod[const2Ftu] 
       (\Nanod[const2Ftu] ), .\Nanod[tvn2Ftu]  (\Nanod[tvn2Ftu] ),
       .\Nanod[clrTpend]  (\Nanod[clrTpend] ), .\Nanod[updTpend] 
       (\Nanod[updTpend] ), .\Nanod[noHighByte]  (\Nanod[noHighByte] ),
       .\Nanod[noLowByte]  (\Nanod[noLowByte] ), .\Nanod[isRmc] 
       (\Nanod[isRmc] ), .\Nanod[busByte]  (\Nanod[busByte] ),
       .\Nanod[isWrite]  (\Nanod[isWrite] ), .\Nanod[waitBusFinish] 
       (\Nanod[waitBusFinish] ), .\Nanod[permStart]  (\Nanod[permStart]
       ), .\Irdecod[inhibitCcr]  (\Irdecod[inhibitCcr] ),
       .\Irdecod[macroTvn]  (\Irdecod[macroTvn] ), .\Irdecod[ftuConst] 
       (\Irdecod[ftuConst] ), .\Irdecod[ryIsAreg]  (\Irdecod[ryIsAreg]
       ), .\Irdecod[rxIsAreg]  (\Irdecod[rxIsAreg] ), .\Irdecod[ry] 
       (\Irdecod[ry] ), .\Irdecod[rx]  (\Irdecod[rx] ),
       .\Irdecod[isMovep]  (\Irdecod[isMovep] ), .\Irdecod[isByte] 
       (\Irdecod[isByte] ), .\Irdecod[movemPreDecr] 
       (\Irdecod[movemPreDecr] ), .\Irdecod[rxIsMovem] 
       (\Irdecod[rxIsMovem] ), .\Irdecod[rxIsUsp]  (\Irdecod[rxIsUsp]
       ), .\Irdecod[ryIsDt]  (\Irdecod[ryIsDt] ), .\Irdecod[rxIsDt] 
       (\Irdecod[rxIsDt] ), .\Irdecod[toCcr]  (\Irdecod[toCcr] ),
       .\Irdecod[implicitSp]  (\Irdecod[implicitSp] ), .\Irdecod[isTas]
        (\Irdecod[isTas] ), .\Irdecod[isPcRel]  (\Irdecod[isPcRel] ),
       .iEdb (iEdb), .aob0 (aob0), .dobIdle (dobIdle), .dobInput
       (dobInput), .Irc (Irc), .dbin (dbin), .oEdb (oEdb));
  fx68k_fx68kAlu alu(.clk (\Clks[clk] ), .pwrUp (\Clks[pwrUp] ), .enT1
       (enT1), .enT3 (enT3), .enT4 (enT4), .ird (Ird), .aluColumn
       (\Nanod[aluColumn] ), .aluDataCtrl (\Nanod[aluDctrl] ),
       .aluAddrCtrl (\Nanod[aluActrl] ), .alueClkEn (alueClkEn),
       .ftu2Ccr (\Nanod[ftu2Ccr] ), .init (\Nanod[aluInit] ), .finish
       (\Nanod[aluFinish] ), .aluIsByte (\Irdecod[isByte] ), .ftu
       (ftu), .alub (alub), .iDataBus (Dbd), .iAddrBus ({Abd[15:3],
       dcrInput[2:0]}), .ze (ze), .alue (alue), .ccr (ccr), .aluOut
       (aluOut));
  fx68k_and_op_1163 g4(.A (rxReg), .Z (n_9));
  fx68k_and_op_1165 g7(.A (ryReg), .Z (n_1344));
  fx68k_bmux_1503 mux_prenLatch_1606_4(.ctl (n_423), .in_0
       (prenLatch[0]), .in_1 (1'b0), .z (n_459));
  fx68k_bmux_1503 mux_prenLatch_1606_129(.ctl (n_424), .in_0
       (prenLatch[1]), .in_1 (1'b0), .z (n_460));
  fx68k_bmux_1503 mux_prenLatch_1606_130(.ctl (n_426), .in_0
       (prenLatch[2]), .in_1 (1'b0), .z (n_461));
  fx68k_bmux_1503 mux_prenLatch_1606_131(.ctl (n_427), .in_0
       (prenLatch[3]), .in_1 (1'b0), .z (n_462));
  fx68k_bmux_1503 mux_prenLatch_1606_132(.ctl (n_428), .in_0
       (prenLatch[4]), .in_1 (1'b0), .z (n_463));
  fx68k_bmux_1503 mux_prenLatch_1606_133(.ctl (n_429), .in_0
       (prenLatch[5]), .in_1 (1'b0), .z (n_464));
  fx68k_bmux_1503 mux_prenLatch_1606_134(.ctl (n_430), .in_0
       (prenLatch[6]), .in_1 (1'b0), .z (n_465));
  fx68k_bmux_1503 mux_prenLatch_1606_135(.ctl (n_431), .in_0
       (prenLatch[7]), .in_1 (1'b0), .z (n_466));
  fx68k_bmux_1503 mux_prenLatch_1606_136(.ctl (n_432), .in_0
       (prenLatch[8]), .in_1 (1'b0), .z (n_467));
  fx68k_bmux_1503 mux_prenLatch_1606_137(.ctl (n_433), .in_0
       (prenLatch[9]), .in_1 (1'b0), .z (n_468));
  fx68k_bmux_1503 mux_prenLatch_1606_138(.ctl (n_434), .in_0
       (prenLatch[10]), .in_1 (1'b0), .z (n_469));
  fx68k_bmux_1503 mux_prenLatch_1606_139(.ctl (n_435), .in_0
       (prenLatch[11]), .in_1 (1'b0), .z (n_470));
  fx68k_bmux_1503 mux_prenLatch_1606_140(.ctl (n_436), .in_0
       (prenLatch[12]), .in_1 (1'b0), .z (n_471));
  fx68k_bmux_1503 mux_prenLatch_1606_141(.ctl (n_437), .in_0
       (prenLatch[13]), .in_1 (1'b0), .z (n_472));
  fx68k_bmux_1503 mux_prenLatch_1606_142(.ctl (n_438), .in_0
       (prenLatch[14]), .in_1 (1'b0), .z (n_473));
  fx68k_bmux_1503 mux_prenLatch_1606_143(.ctl (n_439), .in_0
       (prenLatch[15]), .in_1 (1'b0), .z (n_474));
  fx68k_not_op_1232 g144(.A (prHbit), .Z ({n_478, n_477, n_476,
       n_475}));
  fx68k_add_unsigned_1948 add_1490_27(.A ({Dbh, Dbl}), .B (auInpMux),
       .Z ({n_1265, n_1264, n_1263, n_1262, n_1261, n_1260, n_1259,
       n_1258, n_1257, n_1256, n_1255, n_1254, n_1253, n_1252, n_1251,
       n_1250, n_1249, n_1248, n_1247, n_1246, n_1245, n_1244, n_1243,
       n_1242, n_1241, n_1240, n_1239, n_1238, n_1237, n_1236, n_1235,
       n_1234}));
  fx68k_bmux_1882 mux_prenLatch_1603_12(.ctl (n_456), .in_0 ({n_474,
       n_473, n_472, n_471, n_470, n_469, n_468, n_467, n_466, n_465,
       n_464, n_463, n_462, n_461, n_460, n_459}), .in_1 (dbin), .z
       ({n_6285, n_6284, n_6283, n_6282, n_6281, n_6280, n_6279,
       n_6278, n_6277, n_6276, n_6275, n_6274, n_6273, n_6272, n_6271,
       n_6269}));
  fx68k_bmux_1504 mux_1607_15(.ctl (\Irdecod[movemPreDecr] ), .in_0
       (prHbit), .in_1 ({n_478, n_477, n_476, n_475}), .z ({n_6267,
       n_6266, n_6265, n_6263}));
  fx68k_bmux_1504 mux_rxReg_1241_13(.ctl (\Irdecod[rxIsMovem] ), .in_0
       ({\Irdecod[rxIsAreg] , \Irdecod[rx] }), .in_1 (movemRx), .z
       ({n_486, n_485, n_484, n_483}));
  fx68k_bmux_1504 mux_rxReg_1239_8(.ctl (\Irdecod[implicitSp] ), .in_0
       ({n_486, n_485, n_484, n_483}), .in_1 (4'b1111), .z (rxReg));
  fx68k_mux_1550 mux_rxIsSp_1223_7(.ctl ({\Nanod[ssp] , n_492, n_493,
       n_494, n_495}), .in_0 (1'b1), .in_1 (1'b1), .in_2 (1'b0), .in_3
       (1'b1), .in_4 (1'b0), .z (rxIsSp));
  fx68k_mux_1828 mux_rxMux_1223_7(.ctl ({\Nanod[ssp] , n_492, n_493,
       n_501, n_502, n_503}), .in_0 (5'b10000), .in_1 (5'b01111), .in_2
       (5'b10001), .in_3 (5'b10000), .in_4 (5'b01111), .in_5 ({1'b0,
       rxReg}), .z (rxMux));
  fx68k_bmux_1503 mux_Pcl2Dbl_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_505), .in_1 (1'b0), .z (UNCONNECTED442));
  fx68k_mux_1959 mux_dblIdle_1319_10(.ctl ({rxl2Dbl, ryl2Dbl,
       \Nanod[ftu2Dbl] , \Nanod[au2Db] , \Nanod[atl2Dbl] , Pcl2Dbl,
       n_517}), .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0),
       .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b1), .z (dblIdle));
  fx68k_mux_1550 mux_abdIdle_1338_10(.ctl ({ryl2Abd, rxl2Abd,
       \Nanod[dbin2Abd] , \Nanod[alu2Abd] , n_535}), .in_0 (1'b0),
       .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0), .in_4 (1'b1), .z
       (abdIdle));
  fx68k_bmux_1503 mux_Pcl2Abl_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_537), .in_1 (1'b0), .z (UNCONNECTED443));
  fx68k_mux_1526 mux_ablIdle_1346_10(.ctl ({Pcl2Abl, rxl2Abl, ryl2Abl,
       \Nanod[ftu2Abl] , \Nanod[au2Ab] , \Nanod[aob2Ab] ,
       \Nanod[atl2Abl] , n_551}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b0),
       .in_7 (1'b1), .z (ablIdle));
  fx68k_bmux_1503 mux_dbl2Pcl_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_554), .in_1 (1'b0), .z (UNCONNECTED444));
  fx68k_bmux_1503 mux_abl2Pcl_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_555), .in_1 (1'b0), .z (UNCONNECTED445));
  fx68k_bmux_1882 mux_PcL_1556_8(.ctl (dbl2Pcl), .in_0 (AblOut), .in_1
       (Dbl), .z ({n_587, n_586, n_585, n_584, n_583, n_582, n_581,
       n_580, n_579, n_578, n_577, n_576, n_575, n_574, n_573, n_572}));
  fx68k_bmux_1882 mux_PcL_1553_12(.ctl (n_553), .in_0 ({n_587, n_586,
       n_585, n_584, n_583, n_582, n_581, n_580, n_579, n_578, n_577,
       n_576, n_575, n_574, n_573, n_572}), .in_1 (auReg[15:0]), .z
       ({n_6198, n_6197, n_6196, n_6195, n_6194, n_6193, n_6192,
       n_6191, n_6190, n_6189, n_6188, n_6187, n_6186, n_6185, n_6184,
       n_6182}));
  fx68k_bmux_1967 \mux_regs68L[actualRx]_1348_24 (.ctl (actualRx),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({n_635, n_632, n_629, n_626, n_623, n_620, n_617, n_614, n_611,
       n_608, n_605, n_602, n_599, n_596, n_593, n_590}));
  fx68k_bmux_1967 \mux_regs68L[actualRy]_1349_24 (.ctl (actualRy),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({n_636, n_633, n_630, n_627, n_624, n_621, n_618, n_615, n_612,
       n_609, n_606, n_603, n_600, n_597, n_594, n_591}));
  fx68k_bmux_1882 mux_Atl_1574_8(.ctl (\Nanod[dbl2Atl] ), .in_0
       (AblOut), .in_1 (Dbl), .z ({n_6261, n_6260, n_6259, n_6258,
       n_6257, n_6256, n_6255, n_6254, n_6253, n_6252, n_6251, n_6250,
       n_6249, n_6248, n_6247, n_6245}));
  fx68k_mux_1906 mux_ablMux_1346_10(.ctl ({Pcl2Abl, rxl2Abl, ryl2Abl,
       \Nanod[ftu2Abl] , \Nanod[au2Ab] , \Nanod[aob2Ab] ,
       \Nanod[atl2Abl] }), .in_0 (PcL), .in_1 ({n_635, n_632, n_629,
       n_626, n_623, n_620, n_617, n_614, n_611, n_608, n_605, n_602,
       n_599, n_596, n_593, n_590}), .in_2 ({n_636, n_633, n_630,
       n_627, n_624, n_621, n_618, n_615, n_612, n_609, n_606, n_603,
       n_600, n_597, n_594, n_591}), .in_3 (ftu), .in_4 (auReg[15:0]),
       .in_5 ({eab[15:1], aob0}), .in_6 (Atl), .z (ablMux));
  fx68k_bmux_1503 mux_Pch2Abh_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_639), .in_1 (1'b0), .z (UNCONNECTED446));
  fx68k_bmux_1503 mux_dbh2Pch_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_641), .in_1 (1'b0), .z (UNCONNECTED447));
  fx68k_bmux_1967 \mux_regs68L[actualRy]_1310_24 (.ctl (actualRy),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({\regs68L[actualRy] [15], \regs68L[actualRy] [14],
       \regs68L[actualRy] [13], \regs68L[actualRy] [12],
       \regs68L[actualRy] [11], \regs68L[actualRy] [10],
       \regs68L[actualRy] [9], \regs68L[actualRy] [8],
       \regs68L[actualRy] [7], \regs68L[actualRy] [6],
       \regs68L[actualRy] [5], \regs68L[actualRy] [4],
       \regs68L[actualRy] [3], \regs68L[actualRy] [2],
       \regs68L[actualRy] [1], \regs68L[actualRy] [0]}));
  fx68k_bmux_1967 \mux_regs68L[actualRx]_1311_24 (.ctl (actualRx),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({\regs68L[actualRx] [15], \regs68L[actualRx] [14],
       \regs68L[actualRx] [13], \regs68L[actualRx] [12],
       \regs68L[actualRx] [11], \regs68L[actualRx] [10],
       \regs68L[actualRx] [9], \regs68L[actualRx] [8],
       \regs68L[actualRx] [7], \regs68L[actualRx] [6],
       \regs68L[actualRx] [5], \regs68L[actualRx] [4],
       \regs68L[actualRx] [3], \regs68L[actualRx] [2],
       \regs68L[actualRx] [1], \regs68L[actualRx] [0]}));
  fx68k_bmux_1503 mux_1614_24(.ctl (abdIsByte), .in_0 (Abd[3]), .in_1
       (1'b0), .z (dcrInput[3]));
  fx68k_bmux_1503 mux_Pch2Dbh_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_644), .in_1 (1'b0), .z (UNCONNECTED448));
  fx68k_mux_1707 mux_dbhIdle_1329_10(.ctl ({\Nanod[rxh2dbh] ,
       \Nanod[ryh2dbh] , \Nanod[au2Db] , \Nanod[ath2Dbh] , Pch2Dbh,
       n_653}), .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b0), .in_3 (1'b0),
       .in_4 (1'b0), .in_5 (1'b1), .z (dbhIdle));
  fx68k_mux_1959 mux_abhIdle_1357_10(.ctl ({Pch2Abh, \Nanod[rxh2abh] ,
       \Nanod[ryh2abh] , \Nanod[au2Ab] , \Nanod[aob2Ab] ,
       \Nanod[ath2Abh] , n_666}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b1),
       .z (abhIdle));
  fx68k_bmux_1882 mux_1523_27(.ctl (\Nanod[dbh2ryh] ), .in_0 (Abh),
       .in_1 (Dbh), .z ({n_701, n_699, n_697, n_695, n_693, n_691,
       n_689, n_687, n_685, n_683, n_681, n_679, n_677, n_675, n_673,
       n_671}));
  fx68k_bmux_1882 mux_1521_27(.ctl (\Nanod[dbh2rxh] ), .in_0 (Abh),
       .in_1 (Dbh), .z ({n_702, n_700, n_698, n_696, n_694, n_692,
       n_690, n_688, n_686, n_684, n_682, n_680, n_678, n_676, n_674,
       n_672}));
  fx68k_mux_1995 \mux_regs68H[0]_1523_5 (.ctl ({n_669, n_670}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_718,
       n_717, n_716, n_715, n_714, n_713, n_712, n_711, n_710, n_709,
       n_708, n_707, n_706, n_705, n_704, n_703}));
  fx68k_bmux_1882 \mux_regs68H[0]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_718,
       n_717, n_716, n_715, n_714, n_713, n_712, n_711, n_710, n_709,
       n_708, n_707, n_706, n_705, n_704, n_703}), .z ({n_6175, n_6174,
       n_6173, n_6172, n_6171, n_6170, n_6169, n_6168, n_6167, n_6166,
       n_6165, n_6164, n_6163, n_6162, n_6161, n_6159}));
  fx68k_mux_1995 \mux_regs68H[1]_1523_5 (.ctl ({n_719, n_720}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_736,
       n_735, n_734, n_733, n_732, n_731, n_730, n_729, n_728, n_727,
       n_726, n_725, n_724, n_723, n_722, n_721}));
  fx68k_bmux_1882 \mux_regs68H[1]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_736,
       n_735, n_734, n_733, n_732, n_731, n_730, n_729, n_728, n_727,
       n_726, n_725, n_724, n_723, n_722, n_721}), .z ({n_6151, n_6150,
       n_6149, n_6148, n_6147, n_6146, n_6145, n_6144, n_6143, n_6142,
       n_6141, n_6140, n_6139, n_6138, n_6137, n_6135}));
  fx68k_mux_1995 \mux_regs68H[2]_1523_5 (.ctl ({n_737, n_738}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_754,
       n_753, n_752, n_751, n_750, n_749, n_748, n_747, n_746, n_745,
       n_744, n_743, n_742, n_741, n_740, n_739}));
  fx68k_bmux_1882 \mux_regs68H[2]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_754,
       n_753, n_752, n_751, n_750, n_749, n_748, n_747, n_746, n_745,
       n_744, n_743, n_742, n_741, n_740, n_739}), .z ({n_6127, n_6126,
       n_6125, n_6124, n_6123, n_6122, n_6121, n_6120, n_6119, n_6118,
       n_6117, n_6116, n_6115, n_6114, n_6113, n_6111}));
  fx68k_mux_1995 \mux_regs68H[3]_1523_5 (.ctl ({n_755, n_756}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_772,
       n_771, n_770, n_769, n_768, n_767, n_766, n_765, n_764, n_763,
       n_762, n_761, n_760, n_759, n_758, n_757}));
  fx68k_bmux_1882 \mux_regs68H[3]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_772,
       n_771, n_770, n_769, n_768, n_767, n_766, n_765, n_764, n_763,
       n_762, n_761, n_760, n_759, n_758, n_757}), .z ({n_6103, n_6102,
       n_6101, n_6100, n_6099, n_6098, n_6097, n_6096, n_6095, n_6094,
       n_6093, n_6092, n_6091, n_6090, n_6089, n_6087}));
  fx68k_mux_1995 \mux_regs68H[4]_1523_5 (.ctl ({n_773, n_774}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_790,
       n_789, n_788, n_787, n_786, n_785, n_784, n_783, n_782, n_781,
       n_780, n_779, n_778, n_777, n_776, n_775}));
  fx68k_bmux_1882 \mux_regs68H[4]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_790,
       n_789, n_788, n_787, n_786, n_785, n_784, n_783, n_782, n_781,
       n_780, n_779, n_778, n_777, n_776, n_775}), .z ({n_6079, n_6078,
       n_6077, n_6076, n_6075, n_6074, n_6073, n_6072, n_6071, n_6070,
       n_6069, n_6068, n_6067, n_6066, n_6065, n_6063}));
  fx68k_mux_1995 \mux_regs68H[5]_1523_5 (.ctl ({n_791, n_792}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_808,
       n_807, n_806, n_805, n_804, n_803, n_802, n_801, n_800, n_799,
       n_798, n_797, n_796, n_795, n_794, n_793}));
  fx68k_bmux_1882 \mux_regs68H[5]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_808,
       n_807, n_806, n_805, n_804, n_803, n_802, n_801, n_800, n_799,
       n_798, n_797, n_796, n_795, n_794, n_793}), .z ({n_6055, n_6054,
       n_6053, n_6052, n_6051, n_6050, n_6049, n_6048, n_6047, n_6046,
       n_6045, n_6044, n_6043, n_6042, n_6041, n_6039}));
  fx68k_mux_1995 \mux_regs68H[6]_1523_5 (.ctl ({n_809, n_810}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_826,
       n_825, n_824, n_823, n_822, n_821, n_820, n_819, n_818, n_817,
       n_816, n_815, n_814, n_813, n_812, n_811}));
  fx68k_bmux_1882 \mux_regs68H[6]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_826,
       n_825, n_824, n_823, n_822, n_821, n_820, n_819, n_818, n_817,
       n_816, n_815, n_814, n_813, n_812, n_811}), .z ({n_6031, n_6030,
       n_6029, n_6028, n_6027, n_6026, n_6025, n_6024, n_6023, n_6022,
       n_6021, n_6020, n_6019, n_6018, n_6017, n_6015}));
  fx68k_mux_1995 \mux_regs68H[7]_1523_5 (.ctl ({n_827, n_828}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_844,
       n_843, n_842, n_841, n_840, n_839, n_838, n_837, n_836, n_835,
       n_834, n_833, n_832, n_831, n_830, n_829}));
  fx68k_bmux_1882 \mux_regs68H[7]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_844,
       n_843, n_842, n_841, n_840, n_839, n_838, n_837, n_836, n_835,
       n_834, n_833, n_832, n_831, n_830, n_829}), .z ({n_6007, n_6006,
       n_6005, n_6004, n_6003, n_6002, n_6001, n_6000, n_5999, n_5998,
       n_5997, n_5996, n_5995, n_5994, n_5993, n_5991}));
  fx68k_mux_1995 \mux_regs68H[8]_1523_5 (.ctl ({n_845, n_846}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_862,
       n_861, n_860, n_859, n_858, n_857, n_856, n_855, n_854, n_853,
       n_852, n_851, n_850, n_849, n_848, n_847}));
  fx68k_bmux_1882 \mux_regs68H[8]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_862,
       n_861, n_860, n_859, n_858, n_857, n_856, n_855, n_854, n_853,
       n_852, n_851, n_850, n_849, n_848, n_847}), .z ({n_5983, n_5982,
       n_5981, n_5980, n_5979, n_5978, n_5977, n_5976, n_5975, n_5974,
       n_5973, n_5972, n_5971, n_5970, n_5969, n_5967}));
  fx68k_mux_1995 \mux_regs68H[9]_1523_5 (.ctl ({n_863, n_864}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_880,
       n_879, n_878, n_877, n_876, n_875, n_874, n_873, n_872, n_871,
       n_870, n_869, n_868, n_867, n_866, n_865}));
  fx68k_bmux_1882 \mux_regs68H[9]_1522_22 (.ctl (n_654), .in_0 ({n_702,
       n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686, n_684,
       n_682, n_680, n_678, n_676, n_674, n_672}), .in_1 ({n_880,
       n_879, n_878, n_877, n_876, n_875, n_874, n_873, n_872, n_871,
       n_870, n_869, n_868, n_867, n_866, n_865}), .z ({n_5959, n_5958,
       n_5957, n_5956, n_5955, n_5954, n_5953, n_5952, n_5951, n_5950,
       n_5949, n_5948, n_5947, n_5946, n_5945, n_5943}));
  fx68k_mux_1995 \mux_regs68H[10]_1523_5 (.ctl ({n_881, n_882}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_898,
       n_897, n_896, n_895, n_894, n_893, n_892, n_891, n_890, n_889,
       n_888, n_887, n_886, n_885, n_884, n_883}));
  fx68k_bmux_1882 \mux_regs68H[10]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_898, n_897, n_896, n_895, n_894, n_893, n_892, n_891, n_890,
       n_889, n_888, n_887, n_886, n_885, n_884, n_883}), .z ({n_5935,
       n_5934, n_5933, n_5932, n_5931, n_5930, n_5929, n_5928, n_5927,
       n_5926, n_5925, n_5924, n_5923, n_5922, n_5921, n_5919}));
  fx68k_mux_1995 \mux_regs68H[11]_1523_5 (.ctl ({n_899, n_900}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_916,
       n_915, n_914, n_913, n_912, n_911, n_910, n_909, n_908, n_907,
       n_906, n_905, n_904, n_903, n_902, n_901}));
  fx68k_bmux_1882 \mux_regs68H[11]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_916, n_915, n_914, n_913, n_912, n_911, n_910, n_909, n_908,
       n_907, n_906, n_905, n_904, n_903, n_902, n_901}), .z ({n_5911,
       n_5910, n_5909, n_5908, n_5907, n_5906, n_5905, n_5904, n_5903,
       n_5902, n_5901, n_5900, n_5899, n_5898, n_5897, n_5895}));
  fx68k_mux_1995 \mux_regs68H[12]_1523_5 (.ctl ({n_917, n_918}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_934,
       n_933, n_932, n_931, n_930, n_929, n_928, n_927, n_926, n_925,
       n_924, n_923, n_922, n_921, n_920, n_919}));
  fx68k_bmux_1882 \mux_regs68H[12]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_934, n_933, n_932, n_931, n_930, n_929, n_928, n_927, n_926,
       n_925, n_924, n_923, n_922, n_921, n_920, n_919}), .z ({n_5887,
       n_5886, n_5885, n_5884, n_5883, n_5882, n_5881, n_5880, n_5879,
       n_5878, n_5877, n_5876, n_5875, n_5874, n_5873, n_5871}));
  fx68k_mux_1995 \mux_regs68H[13]_1523_5 (.ctl ({n_935, n_936}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_952,
       n_951, n_950, n_949, n_948, n_947, n_946, n_945, n_944, n_943,
       n_942, n_941, n_940, n_939, n_938, n_937}));
  fx68k_bmux_1882 \mux_regs68H[13]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_952, n_951, n_950, n_949, n_948, n_947, n_946, n_945, n_944,
       n_943, n_942, n_941, n_940, n_939, n_938, n_937}), .z ({n_5863,
       n_5862, n_5861, n_5860, n_5859, n_5858, n_5857, n_5856, n_5855,
       n_5854, n_5853, n_5852, n_5851, n_5850, n_5849, n_5847}));
  fx68k_mux_1995 \mux_regs68H[14]_1523_5 (.ctl ({n_953, n_954}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_970,
       n_969, n_968, n_967, n_966, n_965, n_964, n_963, n_962, n_961,
       n_960, n_959, n_958, n_957, n_956, n_955}));
  fx68k_bmux_1882 \mux_regs68H[14]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_970, n_969, n_968, n_967, n_966, n_965, n_964, n_963, n_962,
       n_961, n_960, n_959, n_958, n_957, n_956, n_955}), .z ({n_5839,
       n_5838, n_5837, n_5836, n_5835, n_5834, n_5833, n_5832, n_5831,
       n_5830, n_5829, n_5828, n_5827, n_5826, n_5825, n_5823}));
  fx68k_mux_1995 \mux_regs68H[15]_1523_5 (.ctl ({n_971, n_972}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_988,
       n_987, n_986, n_985, n_984, n_983, n_982, n_981, n_980, n_979,
       n_978, n_977, n_976, n_975, n_974, n_973}));
  fx68k_bmux_1882 \mux_regs68H[15]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_988, n_987, n_986, n_985, n_984, n_983, n_982, n_981, n_980,
       n_979, n_978, n_977, n_976, n_975, n_974, n_973}), .z ({n_5815,
       n_5814, n_5813, n_5812, n_5811, n_5810, n_5809, n_5808, n_5807,
       n_5806, n_5805, n_5804, n_5803, n_5802, n_5801, n_5799}));
  fx68k_mux_1995 \mux_regs68H[16]_1523_5 (.ctl ({n_989, n_990}), .in_0
       ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687, n_685,
       n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_1006,
       n_1005, n_1004, n_1003, n_1002, n_1001, n_1000, n_999, n_998,
       n_997, n_996, n_995, n_994, n_993, n_992, n_991}));
  fx68k_bmux_1882 \mux_regs68H[16]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_1006, n_1005, n_1004, n_1003, n_1002, n_1001, n_1000, n_999,
       n_998, n_997, n_996, n_995, n_994, n_993, n_992, n_991}), .z
       ({n_5791, n_5790, n_5789, n_5788, n_5787, n_5786, n_5785,
       n_5784, n_5783, n_5782, n_5781, n_5780, n_5779, n_5778, n_5777,
       n_5775}));
  fx68k_mux_1995 \mux_regs68H[17]_1523_5 (.ctl ({n_1007, n_1008}),
       .in_0 ({n_701, n_699, n_697, n_695, n_693, n_691, n_689, n_687,
       n_685, n_683, n_681, n_679, n_677, n_675, n_673, n_671}), .in_1
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .z ({n_1024,
       n_1023, n_1022, n_1021, n_1020, n_1019, n_1018, n_1017, n_1016,
       n_1015, n_1014, n_1013, n_1012, n_1011, n_1010, n_1009}));
  fx68k_bmux_1882 \mux_regs68H[17]_1522_22 (.ctl (n_654), .in_0
       ({n_702, n_700, n_698, n_696, n_694, n_692, n_690, n_688, n_686,
       n_684, n_682, n_680, n_678, n_676, n_674, n_672}), .in_1
       ({n_1024, n_1023, n_1022, n_1021, n_1020, n_1019, n_1018,
       n_1017, n_1016, n_1015, n_1014, n_1013, n_1012, n_1011, n_1010,
       n_1009}), .z ({n_5767, n_5766, n_5765, n_5764, n_5763, n_5762,
       n_5761, n_5760, n_5759, n_5758, n_5757, n_5756, n_5755, n_5754,
       n_5753, n_5751}));
  fx68k_bmux_1967 \mux_regs68H[actualRx]_1330_29 (.ctl (actualRx),
       .in_0 ({\regs68H[0] [15], \regs68H[0] [14], \regs68H[0] [13],
       \regs68H[0] [12], \regs68H[0] [11], \regs68H[0] [10],
       \regs68H[0] [9], \regs68H[0] [8], \regs68H[0] [7],
       \regs68H[0] [6], \regs68H[0] [5], \regs68H[0] [4],
       \regs68H[0] [3], \regs68H[0] [2], \regs68H[0] [1],
       \regs68H[0] [0]}), .in_1 ({\regs68H[1] [15], \regs68H[1] [14],
       \regs68H[1] [13], \regs68H[1] [12], \regs68H[1] [11],
       \regs68H[1] [10], \regs68H[1] [9], \regs68H[1] [8],
       \regs68H[1] [7], \regs68H[1] [6], \regs68H[1] [5],
       \regs68H[1] [4], \regs68H[1] [3], \regs68H[1] [2],
       \regs68H[1] [1], \regs68H[1] [0]}), .in_2 ({\regs68H[2] [15],
       \regs68H[2] [14], \regs68H[2] [13], \regs68H[2] [12],
       \regs68H[2] [11], \regs68H[2] [10], \regs68H[2] [9],
       \regs68H[2] [8], \regs68H[2] [7], \regs68H[2] [6],
       \regs68H[2] [5], \regs68H[2] [4], \regs68H[2] [3],
       \regs68H[2] [2], \regs68H[2] [1], \regs68H[2] [0]}), .in_3
       ({\regs68H[3] [15], \regs68H[3] [14], \regs68H[3] [13],
       \regs68H[3] [12], \regs68H[3] [11], \regs68H[3] [10],
       \regs68H[3] [9], \regs68H[3] [8], \regs68H[3] [7],
       \regs68H[3] [6], \regs68H[3] [5], \regs68H[3] [4],
       \regs68H[3] [3], \regs68H[3] [2], \regs68H[3] [1],
       \regs68H[3] [0]}), .in_4 ({\regs68H[4] [15], \regs68H[4] [14],
       \regs68H[4] [13], \regs68H[4] [12], \regs68H[4] [11],
       \regs68H[4] [10], \regs68H[4] [9], \regs68H[4] [8],
       \regs68H[4] [7], \regs68H[4] [6], \regs68H[4] [5],
       \regs68H[4] [4], \regs68H[4] [3], \regs68H[4] [2],
       \regs68H[4] [1], \regs68H[4] [0]}), .in_5 ({\regs68H[5] [15],
       \regs68H[5] [14], \regs68H[5] [13], \regs68H[5] [12],
       \regs68H[5] [11], \regs68H[5] [10], \regs68H[5] [9],
       \regs68H[5] [8], \regs68H[5] [7], \regs68H[5] [6],
       \regs68H[5] [5], \regs68H[5] [4], \regs68H[5] [3],
       \regs68H[5] [2], \regs68H[5] [1], \regs68H[5] [0]}), .in_6
       ({\regs68H[6] [15], \regs68H[6] [14], \regs68H[6] [13],
       \regs68H[6] [12], \regs68H[6] [11], \regs68H[6] [10],
       \regs68H[6] [9], \regs68H[6] [8], \regs68H[6] [7],
       \regs68H[6] [6], \regs68H[6] [5], \regs68H[6] [4],
       \regs68H[6] [3], \regs68H[6] [2], \regs68H[6] [1],
       \regs68H[6] [0]}), .in_7 ({\regs68H[7] [15], \regs68H[7] [14],
       \regs68H[7] [13], \regs68H[7] [12], \regs68H[7] [11],
       \regs68H[7] [10], \regs68H[7] [9], \regs68H[7] [8],
       \regs68H[7] [7], \regs68H[7] [6], \regs68H[7] [5],
       \regs68H[7] [4], \regs68H[7] [3], \regs68H[7] [2],
       \regs68H[7] [1], \regs68H[7] [0]}), .in_8 ({\regs68H[8] [15],
       \regs68H[8] [14], \regs68H[8] [13], \regs68H[8] [12],
       \regs68H[8] [11], \regs68H[8] [10], \regs68H[8] [9],
       \regs68H[8] [8], \regs68H[8] [7], \regs68H[8] [6],
       \regs68H[8] [5], \regs68H[8] [4], \regs68H[8] [3],
       \regs68H[8] [2], \regs68H[8] [1], \regs68H[8] [0]}), .in_9
       ({\regs68H[9] [15], \regs68H[9] [14], \regs68H[9] [13],
       \regs68H[9] [12], \regs68H[9] [11], \regs68H[9] [10],
       \regs68H[9] [9], \regs68H[9] [8], \regs68H[9] [7],
       \regs68H[9] [6], \regs68H[9] [5], \regs68H[9] [4],
       \regs68H[9] [3], \regs68H[9] [2], \regs68H[9] [1],
       \regs68H[9] [0]}), .in_10 ({\regs68H[10] [15], \regs68H[10]
       [14], \regs68H[10] [13], \regs68H[10] [12], \regs68H[10] [11],
       \regs68H[10] [10], \regs68H[10] [9], \regs68H[10] [8],
       \regs68H[10] [7], \regs68H[10] [6], \regs68H[10] [5],
       \regs68H[10] [4], \regs68H[10] [3], \regs68H[10] [2],
       \regs68H[10] [1], \regs68H[10] [0]}), .in_11 ({\regs68H[11]
       [15], \regs68H[11] [14], \regs68H[11] [13], \regs68H[11] [12],
       \regs68H[11] [11], \regs68H[11] [10], \regs68H[11] [9],
       \regs68H[11] [8], \regs68H[11] [7], \regs68H[11] [6],
       \regs68H[11] [5], \regs68H[11] [4], \regs68H[11] [3],
       \regs68H[11] [2], \regs68H[11] [1], \regs68H[11] [0]}), .in_12
       ({\regs68H[12] [15], \regs68H[12] [14], \regs68H[12] [13],
       \regs68H[12] [12], \regs68H[12] [11], \regs68H[12] [10],
       \regs68H[12] [9], \regs68H[12] [8], \regs68H[12] [7],
       \regs68H[12] [6], \regs68H[12] [5], \regs68H[12] [4],
       \regs68H[12] [3], \regs68H[12] [2], \regs68H[12] [1],
       \regs68H[12] [0]}), .in_13 ({\regs68H[13] [15], \regs68H[13]
       [14], \regs68H[13] [13], \regs68H[13] [12], \regs68H[13] [11],
       \regs68H[13] [10], \regs68H[13] [9], \regs68H[13] [8],
       \regs68H[13] [7], \regs68H[13] [6], \regs68H[13] [5],
       \regs68H[13] [4], \regs68H[13] [3], \regs68H[13] [2],
       \regs68H[13] [1], \regs68H[13] [0]}), .in_14 ({\regs68H[14]
       [15], \regs68H[14] [14], \regs68H[14] [13], \regs68H[14] [12],
       \regs68H[14] [11], \regs68H[14] [10], \regs68H[14] [9],
       \regs68H[14] [8], \regs68H[14] [7], \regs68H[14] [6],
       \regs68H[14] [5], \regs68H[14] [4], \regs68H[14] [3],
       \regs68H[14] [2], \regs68H[14] [1], \regs68H[14] [0]}), .in_15
       ({\regs68H[15] [15], \regs68H[15] [14], \regs68H[15] [13],
       \regs68H[15] [12], \regs68H[15] [11], \regs68H[15] [10],
       \regs68H[15] [9], \regs68H[15] [8], \regs68H[15] [7],
       \regs68H[15] [6], \regs68H[15] [5], \regs68H[15] [4],
       \regs68H[15] [3], \regs68H[15] [2], \regs68H[15] [1],
       \regs68H[15] [0]}), .in_16 ({\regs68H[16] [15], \regs68H[16]
       [14], \regs68H[16] [13], \regs68H[16] [12], \regs68H[16] [11],
       \regs68H[16] [10], \regs68H[16] [9], \regs68H[16] [8],
       \regs68H[16] [7], \regs68H[16] [6], \regs68H[16] [5],
       \regs68H[16] [4], \regs68H[16] [3], \regs68H[16] [2],
       \regs68H[16] [1], \regs68H[16] [0]}), .in_17 ({\regs68H[17]
       [15], \regs68H[17] [14], \regs68H[17] [13], \regs68H[17] [12],
       \regs68H[17] [11], \regs68H[17] [10], \regs68H[17] [9],
       \regs68H[17] [8], \regs68H[17] [7], \regs68H[17] [6],
       \regs68H[17] [5], \regs68H[17] [4], \regs68H[17] [3],
       \regs68H[17] [2], \regs68H[17] [1], \regs68H[17] [0]}), .z
       ({\regs68H[actualRx] [15], \regs68H[actualRx] [14],
       \regs68H[actualRx] [13], \regs68H[actualRx] [12],
       \regs68H[actualRx] [11], \regs68H[actualRx] [10],
       \regs68H[actualRx] [9], \regs68H[actualRx] [8],
       \regs68H[actualRx] [7], \regs68H[actualRx] [6],
       \regs68H[actualRx] [5], \regs68H[actualRx] [4],
       \regs68H[actualRx] [3], \regs68H[actualRx] [2],
       \regs68H[actualRx] [1], \regs68H[actualRx] [0]}));
  fx68k_bmux_1967 \mux_regs68H[actualRy]_1331_29 (.ctl (actualRy),
       .in_0 ({\regs68H[0] [15], \regs68H[0] [14], \regs68H[0] [13],
       \regs68H[0] [12], \regs68H[0] [11], \regs68H[0] [10],
       \regs68H[0] [9], \regs68H[0] [8], \regs68H[0] [7],
       \regs68H[0] [6], \regs68H[0] [5], \regs68H[0] [4],
       \regs68H[0] [3], \regs68H[0] [2], \regs68H[0] [1],
       \regs68H[0] [0]}), .in_1 ({\regs68H[1] [15], \regs68H[1] [14],
       \regs68H[1] [13], \regs68H[1] [12], \regs68H[1] [11],
       \regs68H[1] [10], \regs68H[1] [9], \regs68H[1] [8],
       \regs68H[1] [7], \regs68H[1] [6], \regs68H[1] [5],
       \regs68H[1] [4], \regs68H[1] [3], \regs68H[1] [2],
       \regs68H[1] [1], \regs68H[1] [0]}), .in_2 ({\regs68H[2] [15],
       \regs68H[2] [14], \regs68H[2] [13], \regs68H[2] [12],
       \regs68H[2] [11], \regs68H[2] [10], \regs68H[2] [9],
       \regs68H[2] [8], \regs68H[2] [7], \regs68H[2] [6],
       \regs68H[2] [5], \regs68H[2] [4], \regs68H[2] [3],
       \regs68H[2] [2], \regs68H[2] [1], \regs68H[2] [0]}), .in_3
       ({\regs68H[3] [15], \regs68H[3] [14], \regs68H[3] [13],
       \regs68H[3] [12], \regs68H[3] [11], \regs68H[3] [10],
       \regs68H[3] [9], \regs68H[3] [8], \regs68H[3] [7],
       \regs68H[3] [6], \regs68H[3] [5], \regs68H[3] [4],
       \regs68H[3] [3], \regs68H[3] [2], \regs68H[3] [1],
       \regs68H[3] [0]}), .in_4 ({\regs68H[4] [15], \regs68H[4] [14],
       \regs68H[4] [13], \regs68H[4] [12], \regs68H[4] [11],
       \regs68H[4] [10], \regs68H[4] [9], \regs68H[4] [8],
       \regs68H[4] [7], \regs68H[4] [6], \regs68H[4] [5],
       \regs68H[4] [4], \regs68H[4] [3], \regs68H[4] [2],
       \regs68H[4] [1], \regs68H[4] [0]}), .in_5 ({\regs68H[5] [15],
       \regs68H[5] [14], \regs68H[5] [13], \regs68H[5] [12],
       \regs68H[5] [11], \regs68H[5] [10], \regs68H[5] [9],
       \regs68H[5] [8], \regs68H[5] [7], \regs68H[5] [6],
       \regs68H[5] [5], \regs68H[5] [4], \regs68H[5] [3],
       \regs68H[5] [2], \regs68H[5] [1], \regs68H[5] [0]}), .in_6
       ({\regs68H[6] [15], \regs68H[6] [14], \regs68H[6] [13],
       \regs68H[6] [12], \regs68H[6] [11], \regs68H[6] [10],
       \regs68H[6] [9], \regs68H[6] [8], \regs68H[6] [7],
       \regs68H[6] [6], \regs68H[6] [5], \regs68H[6] [4],
       \regs68H[6] [3], \regs68H[6] [2], \regs68H[6] [1],
       \regs68H[6] [0]}), .in_7 ({\regs68H[7] [15], \regs68H[7] [14],
       \regs68H[7] [13], \regs68H[7] [12], \regs68H[7] [11],
       \regs68H[7] [10], \regs68H[7] [9], \regs68H[7] [8],
       \regs68H[7] [7], \regs68H[7] [6], \regs68H[7] [5],
       \regs68H[7] [4], \regs68H[7] [3], \regs68H[7] [2],
       \regs68H[7] [1], \regs68H[7] [0]}), .in_8 ({\regs68H[8] [15],
       \regs68H[8] [14], \regs68H[8] [13], \regs68H[8] [12],
       \regs68H[8] [11], \regs68H[8] [10], \regs68H[8] [9],
       \regs68H[8] [8], \regs68H[8] [7], \regs68H[8] [6],
       \regs68H[8] [5], \regs68H[8] [4], \regs68H[8] [3],
       \regs68H[8] [2], \regs68H[8] [1], \regs68H[8] [0]}), .in_9
       ({\regs68H[9] [15], \regs68H[9] [14], \regs68H[9] [13],
       \regs68H[9] [12], \regs68H[9] [11], \regs68H[9] [10],
       \regs68H[9] [9], \regs68H[9] [8], \regs68H[9] [7],
       \regs68H[9] [6], \regs68H[9] [5], \regs68H[9] [4],
       \regs68H[9] [3], \regs68H[9] [2], \regs68H[9] [1],
       \regs68H[9] [0]}), .in_10 ({\regs68H[10] [15], \regs68H[10]
       [14], \regs68H[10] [13], \regs68H[10] [12], \regs68H[10] [11],
       \regs68H[10] [10], \regs68H[10] [9], \regs68H[10] [8],
       \regs68H[10] [7], \regs68H[10] [6], \regs68H[10] [5],
       \regs68H[10] [4], \regs68H[10] [3], \regs68H[10] [2],
       \regs68H[10] [1], \regs68H[10] [0]}), .in_11 ({\regs68H[11]
       [15], \regs68H[11] [14], \regs68H[11] [13], \regs68H[11] [12],
       \regs68H[11] [11], \regs68H[11] [10], \regs68H[11] [9],
       \regs68H[11] [8], \regs68H[11] [7], \regs68H[11] [6],
       \regs68H[11] [5], \regs68H[11] [4], \regs68H[11] [3],
       \regs68H[11] [2], \regs68H[11] [1], \regs68H[11] [0]}), .in_12
       ({\regs68H[12] [15], \regs68H[12] [14], \regs68H[12] [13],
       \regs68H[12] [12], \regs68H[12] [11], \regs68H[12] [10],
       \regs68H[12] [9], \regs68H[12] [8], \regs68H[12] [7],
       \regs68H[12] [6], \regs68H[12] [5], \regs68H[12] [4],
       \regs68H[12] [3], \regs68H[12] [2], \regs68H[12] [1],
       \regs68H[12] [0]}), .in_13 ({\regs68H[13] [15], \regs68H[13]
       [14], \regs68H[13] [13], \regs68H[13] [12], \regs68H[13] [11],
       \regs68H[13] [10], \regs68H[13] [9], \regs68H[13] [8],
       \regs68H[13] [7], \regs68H[13] [6], \regs68H[13] [5],
       \regs68H[13] [4], \regs68H[13] [3], \regs68H[13] [2],
       \regs68H[13] [1], \regs68H[13] [0]}), .in_14 ({\regs68H[14]
       [15], \regs68H[14] [14], \regs68H[14] [13], \regs68H[14] [12],
       \regs68H[14] [11], \regs68H[14] [10], \regs68H[14] [9],
       \regs68H[14] [8], \regs68H[14] [7], \regs68H[14] [6],
       \regs68H[14] [5], \regs68H[14] [4], \regs68H[14] [3],
       \regs68H[14] [2], \regs68H[14] [1], \regs68H[14] [0]}), .in_15
       ({\regs68H[15] [15], \regs68H[15] [14], \regs68H[15] [13],
       \regs68H[15] [12], \regs68H[15] [11], \regs68H[15] [10],
       \regs68H[15] [9], \regs68H[15] [8], \regs68H[15] [7],
       \regs68H[15] [6], \regs68H[15] [5], \regs68H[15] [4],
       \regs68H[15] [3], \regs68H[15] [2], \regs68H[15] [1],
       \regs68H[15] [0]}), .in_16 ({\regs68H[16] [15], \regs68H[16]
       [14], \regs68H[16] [13], \regs68H[16] [12], \regs68H[16] [11],
       \regs68H[16] [10], \regs68H[16] [9], \regs68H[16] [8],
       \regs68H[16] [7], \regs68H[16] [6], \regs68H[16] [5],
       \regs68H[16] [4], \regs68H[16] [3], \regs68H[16] [2],
       \regs68H[16] [1], \regs68H[16] [0]}), .in_17 ({\regs68H[17]
       [15], \regs68H[17] [14], \regs68H[17] [13], \regs68H[17] [12],
       \regs68H[17] [11], \regs68H[17] [10], \regs68H[17] [9],
       \regs68H[17] [8], \regs68H[17] [7], \regs68H[17] [6],
       \regs68H[17] [5], \regs68H[17] [4], \regs68H[17] [3],
       \regs68H[17] [2], \regs68H[17] [1], \regs68H[17] [0]}), .z
       ({\regs68H[actualRy] [15], \regs68H[actualRy] [14],
       \regs68H[actualRy] [13], \regs68H[actualRy] [12],
       \regs68H[actualRy] [11], \regs68H[actualRy] [10],
       \regs68H[actualRy] [9], \regs68H[actualRy] [8],
       \regs68H[actualRy] [7], \regs68H[actualRy] [6],
       \regs68H[actualRy] [5], \regs68H[actualRy] [4],
       \regs68H[actualRy] [3], \regs68H[actualRy] [2],
       \regs68H[actualRy] [1], \regs68H[actualRy] [0]}));
  fx68k_bmux_1882 mux_Ath_1582_8(.ctl (\Nanod[abh2Ath] ), .in_0 (Dbh),
       .in_1 (Abh), .z ({n_6241, n_6240, n_6239, n_6238, n_6237,
       n_6236, n_6235, n_6234, n_6233, n_6232, n_6231, n_6230, n_6229,
       n_6228, n_6227, n_6225}));
  fx68k_mux_2286 mux_dbhMux_1329_10(.ctl ({\Nanod[rxh2dbh] ,
       \Nanod[ryh2dbh] , \Nanod[au2Db] , \Nanod[ath2Dbh] , Pch2Dbh}),
       .in_0 ({\regs68H[actualRx] [15], \regs68H[actualRx] [14],
       \regs68H[actualRx] [13], \regs68H[actualRx] [12],
       \regs68H[actualRx] [11], \regs68H[actualRx] [10],
       \regs68H[actualRx] [9], \regs68H[actualRx] [8],
       \regs68H[actualRx] [7], \regs68H[actualRx] [6],
       \regs68H[actualRx] [5], \regs68H[actualRx] [4],
       \regs68H[actualRx] [3], \regs68H[actualRx] [2],
       \regs68H[actualRx] [1], \regs68H[actualRx] [0]}), .in_1
       ({\regs68H[actualRy] [15], \regs68H[actualRy] [14],
       \regs68H[actualRy] [13], \regs68H[actualRy] [12],
       \regs68H[actualRy] [11], \regs68H[actualRy] [10],
       \regs68H[actualRy] [9], \regs68H[actualRy] [8],
       \regs68H[actualRy] [7], \regs68H[actualRy] [6],
       \regs68H[actualRy] [5], \regs68H[actualRy] [4],
       \regs68H[actualRy] [3], \regs68H[actualRy] [2],
       \regs68H[actualRy] [1], \regs68H[actualRy] [0]}), .in_2
       (auReg[31:16]), .in_3 (Ath), .in_4 (PcH), .z (dbhMux));
  fx68k_bmux_1503 mux_abh2Pch_1532_7(.ctl (\Clks[extReset] ), .in_0
       (n_1027), .in_1 (1'b0), .z (UNCONNECTED449));
  fx68k_bmux_1882 mux_PcH_1566_8(.ctl (dbh2Pch), .in_0 (Abh), .in_1
       (Dbh), .z ({n_1043, n_1042, n_1041, n_1040, n_1039, n_1038,
       n_1037, n_1036, n_1035, n_1034, n_1033, n_1032, n_1031, n_1030,
       n_1029, n_1028}));
  fx68k_bmux_1882 mux_PcH_1563_12(.ctl (n_553), .in_0 ({n_1043, n_1042,
       n_1041, n_1040, n_1039, n_1038, n_1037, n_1036, n_1035, n_1034,
       n_1033, n_1032, n_1031, n_1030, n_1029, n_1028}), .in_1
       (auReg[31:16]), .z ({n_6221, n_6220, n_6219, n_6218, n_6217,
       n_6216, n_6215, n_6214, n_6213, n_6212, n_6211, n_6210, n_6209,
       n_6208, n_6207, n_6205}));
  fx68k_bmux_1967 \mux_regs68H[actualRx]_1359_29 (.ctl (actualRx),
       .in_0 ({\regs68H[0] [15], \regs68H[0] [14], \regs68H[0] [13],
       \regs68H[0] [12], \regs68H[0] [11], \regs68H[0] [10],
       \regs68H[0] [9], \regs68H[0] [8], \regs68H[0] [7],
       \regs68H[0] [6], \regs68H[0] [5], \regs68H[0] [4],
       \regs68H[0] [3], \regs68H[0] [2], \regs68H[0] [1],
       \regs68H[0] [0]}), .in_1 ({\regs68H[1] [15], \regs68H[1] [14],
       \regs68H[1] [13], \regs68H[1] [12], \regs68H[1] [11],
       \regs68H[1] [10], \regs68H[1] [9], \regs68H[1] [8],
       \regs68H[1] [7], \regs68H[1] [6], \regs68H[1] [5],
       \regs68H[1] [4], \regs68H[1] [3], \regs68H[1] [2],
       \regs68H[1] [1], \regs68H[1] [0]}), .in_2 ({\regs68H[2] [15],
       \regs68H[2] [14], \regs68H[2] [13], \regs68H[2] [12],
       \regs68H[2] [11], \regs68H[2] [10], \regs68H[2] [9],
       \regs68H[2] [8], \regs68H[2] [7], \regs68H[2] [6],
       \regs68H[2] [5], \regs68H[2] [4], \regs68H[2] [3],
       \regs68H[2] [2], \regs68H[2] [1], \regs68H[2] [0]}), .in_3
       ({\regs68H[3] [15], \regs68H[3] [14], \regs68H[3] [13],
       \regs68H[3] [12], \regs68H[3] [11], \regs68H[3] [10],
       \regs68H[3] [9], \regs68H[3] [8], \regs68H[3] [7],
       \regs68H[3] [6], \regs68H[3] [5], \regs68H[3] [4],
       \regs68H[3] [3], \regs68H[3] [2], \regs68H[3] [1],
       \regs68H[3] [0]}), .in_4 ({\regs68H[4] [15], \regs68H[4] [14],
       \regs68H[4] [13], \regs68H[4] [12], \regs68H[4] [11],
       \regs68H[4] [10], \regs68H[4] [9], \regs68H[4] [8],
       \regs68H[4] [7], \regs68H[4] [6], \regs68H[4] [5],
       \regs68H[4] [4], \regs68H[4] [3], \regs68H[4] [2],
       \regs68H[4] [1], \regs68H[4] [0]}), .in_5 ({\regs68H[5] [15],
       \regs68H[5] [14], \regs68H[5] [13], \regs68H[5] [12],
       \regs68H[5] [11], \regs68H[5] [10], \regs68H[5] [9],
       \regs68H[5] [8], \regs68H[5] [7], \regs68H[5] [6],
       \regs68H[5] [5], \regs68H[5] [4], \regs68H[5] [3],
       \regs68H[5] [2], \regs68H[5] [1], \regs68H[5] [0]}), .in_6
       ({\regs68H[6] [15], \regs68H[6] [14], \regs68H[6] [13],
       \regs68H[6] [12], \regs68H[6] [11], \regs68H[6] [10],
       \regs68H[6] [9], \regs68H[6] [8], \regs68H[6] [7],
       \regs68H[6] [6], \regs68H[6] [5], \regs68H[6] [4],
       \regs68H[6] [3], \regs68H[6] [2], \regs68H[6] [1],
       \regs68H[6] [0]}), .in_7 ({\regs68H[7] [15], \regs68H[7] [14],
       \regs68H[7] [13], \regs68H[7] [12], \regs68H[7] [11],
       \regs68H[7] [10], \regs68H[7] [9], \regs68H[7] [8],
       \regs68H[7] [7], \regs68H[7] [6], \regs68H[7] [5],
       \regs68H[7] [4], \regs68H[7] [3], \regs68H[7] [2],
       \regs68H[7] [1], \regs68H[7] [0]}), .in_8 ({\regs68H[8] [15],
       \regs68H[8] [14], \regs68H[8] [13], \regs68H[8] [12],
       \regs68H[8] [11], \regs68H[8] [10], \regs68H[8] [9],
       \regs68H[8] [8], \regs68H[8] [7], \regs68H[8] [6],
       \regs68H[8] [5], \regs68H[8] [4], \regs68H[8] [3],
       \regs68H[8] [2], \regs68H[8] [1], \regs68H[8] [0]}), .in_9
       ({\regs68H[9] [15], \regs68H[9] [14], \regs68H[9] [13],
       \regs68H[9] [12], \regs68H[9] [11], \regs68H[9] [10],
       \regs68H[9] [9], \regs68H[9] [8], \regs68H[9] [7],
       \regs68H[9] [6], \regs68H[9] [5], \regs68H[9] [4],
       \regs68H[9] [3], \regs68H[9] [2], \regs68H[9] [1],
       \regs68H[9] [0]}), .in_10 ({\regs68H[10] [15], \regs68H[10]
       [14], \regs68H[10] [13], \regs68H[10] [12], \regs68H[10] [11],
       \regs68H[10] [10], \regs68H[10] [9], \regs68H[10] [8],
       \regs68H[10] [7], \regs68H[10] [6], \regs68H[10] [5],
       \regs68H[10] [4], \regs68H[10] [3], \regs68H[10] [2],
       \regs68H[10] [1], \regs68H[10] [0]}), .in_11 ({\regs68H[11]
       [15], \regs68H[11] [14], \regs68H[11] [13], \regs68H[11] [12],
       \regs68H[11] [11], \regs68H[11] [10], \regs68H[11] [9],
       \regs68H[11] [8], \regs68H[11] [7], \regs68H[11] [6],
       \regs68H[11] [5], \regs68H[11] [4], \regs68H[11] [3],
       \regs68H[11] [2], \regs68H[11] [1], \regs68H[11] [0]}), .in_12
       ({\regs68H[12] [15], \regs68H[12] [14], \regs68H[12] [13],
       \regs68H[12] [12], \regs68H[12] [11], \regs68H[12] [10],
       \regs68H[12] [9], \regs68H[12] [8], \regs68H[12] [7],
       \regs68H[12] [6], \regs68H[12] [5], \regs68H[12] [4],
       \regs68H[12] [3], \regs68H[12] [2], \regs68H[12] [1],
       \regs68H[12] [0]}), .in_13 ({\regs68H[13] [15], \regs68H[13]
       [14], \regs68H[13] [13], \regs68H[13] [12], \regs68H[13] [11],
       \regs68H[13] [10], \regs68H[13] [9], \regs68H[13] [8],
       \regs68H[13] [7], \regs68H[13] [6], \regs68H[13] [5],
       \regs68H[13] [4], \regs68H[13] [3], \regs68H[13] [2],
       \regs68H[13] [1], \regs68H[13] [0]}), .in_14 ({\regs68H[14]
       [15], \regs68H[14] [14], \regs68H[14] [13], \regs68H[14] [12],
       \regs68H[14] [11], \regs68H[14] [10], \regs68H[14] [9],
       \regs68H[14] [8], \regs68H[14] [7], \regs68H[14] [6],
       \regs68H[14] [5], \regs68H[14] [4], \regs68H[14] [3],
       \regs68H[14] [2], \regs68H[14] [1], \regs68H[14] [0]}), .in_15
       ({\regs68H[15] [15], \regs68H[15] [14], \regs68H[15] [13],
       \regs68H[15] [12], \regs68H[15] [11], \regs68H[15] [10],
       \regs68H[15] [9], \regs68H[15] [8], \regs68H[15] [7],
       \regs68H[15] [6], \regs68H[15] [5], \regs68H[15] [4],
       \regs68H[15] [3], \regs68H[15] [2], \regs68H[15] [1],
       \regs68H[15] [0]}), .in_16 ({\regs68H[16] [15], \regs68H[16]
       [14], \regs68H[16] [13], \regs68H[16] [12], \regs68H[16] [11],
       \regs68H[16] [10], \regs68H[16] [9], \regs68H[16] [8],
       \regs68H[16] [7], \regs68H[16] [6], \regs68H[16] [5],
       \regs68H[16] [4], \regs68H[16] [3], \regs68H[16] [2],
       \regs68H[16] [1], \regs68H[16] [0]}), .in_17 ({\regs68H[17]
       [15], \regs68H[17] [14], \regs68H[17] [13], \regs68H[17] [12],
       \regs68H[17] [11], \regs68H[17] [10], \regs68H[17] [9],
       \regs68H[17] [8], \regs68H[17] [7], \regs68H[17] [6],
       \regs68H[17] [5], \regs68H[17] [4], \regs68H[17] [3],
       \regs68H[17] [2], \regs68H[17] [1], \regs68H[17] [0]}), .z
       ({n_1074, n_1072, n_1070, n_1068, n_1066, n_1064, n_1062,
       n_1060, n_1058, n_1056, n_1054, n_1052, n_1050, n_1048, n_1046,
       n_1044}));
  fx68k_bmux_1967 \mux_regs68H[actualRy]_1360_29 (.ctl (actualRy),
       .in_0 ({\regs68H[0] [15], \regs68H[0] [14], \regs68H[0] [13],
       \regs68H[0] [12], \regs68H[0] [11], \regs68H[0] [10],
       \regs68H[0] [9], \regs68H[0] [8], \regs68H[0] [7],
       \regs68H[0] [6], \regs68H[0] [5], \regs68H[0] [4],
       \regs68H[0] [3], \regs68H[0] [2], \regs68H[0] [1],
       \regs68H[0] [0]}), .in_1 ({\regs68H[1] [15], \regs68H[1] [14],
       \regs68H[1] [13], \regs68H[1] [12], \regs68H[1] [11],
       \regs68H[1] [10], \regs68H[1] [9], \regs68H[1] [8],
       \regs68H[1] [7], \regs68H[1] [6], \regs68H[1] [5],
       \regs68H[1] [4], \regs68H[1] [3], \regs68H[1] [2],
       \regs68H[1] [1], \regs68H[1] [0]}), .in_2 ({\regs68H[2] [15],
       \regs68H[2] [14], \regs68H[2] [13], \regs68H[2] [12],
       \regs68H[2] [11], \regs68H[2] [10], \regs68H[2] [9],
       \regs68H[2] [8], \regs68H[2] [7], \regs68H[2] [6],
       \regs68H[2] [5], \regs68H[2] [4], \regs68H[2] [3],
       \regs68H[2] [2], \regs68H[2] [1], \regs68H[2] [0]}), .in_3
       ({\regs68H[3] [15], \regs68H[3] [14], \regs68H[3] [13],
       \regs68H[3] [12], \regs68H[3] [11], \regs68H[3] [10],
       \regs68H[3] [9], \regs68H[3] [8], \regs68H[3] [7],
       \regs68H[3] [6], \regs68H[3] [5], \regs68H[3] [4],
       \regs68H[3] [3], \regs68H[3] [2], \regs68H[3] [1],
       \regs68H[3] [0]}), .in_4 ({\regs68H[4] [15], \regs68H[4] [14],
       \regs68H[4] [13], \regs68H[4] [12], \regs68H[4] [11],
       \regs68H[4] [10], \regs68H[4] [9], \regs68H[4] [8],
       \regs68H[4] [7], \regs68H[4] [6], \regs68H[4] [5],
       \regs68H[4] [4], \regs68H[4] [3], \regs68H[4] [2],
       \regs68H[4] [1], \regs68H[4] [0]}), .in_5 ({\regs68H[5] [15],
       \regs68H[5] [14], \regs68H[5] [13], \regs68H[5] [12],
       \regs68H[5] [11], \regs68H[5] [10], \regs68H[5] [9],
       \regs68H[5] [8], \regs68H[5] [7], \regs68H[5] [6],
       \regs68H[5] [5], \regs68H[5] [4], \regs68H[5] [3],
       \regs68H[5] [2], \regs68H[5] [1], \regs68H[5] [0]}), .in_6
       ({\regs68H[6] [15], \regs68H[6] [14], \regs68H[6] [13],
       \regs68H[6] [12], \regs68H[6] [11], \regs68H[6] [10],
       \regs68H[6] [9], \regs68H[6] [8], \regs68H[6] [7],
       \regs68H[6] [6], \regs68H[6] [5], \regs68H[6] [4],
       \regs68H[6] [3], \regs68H[6] [2], \regs68H[6] [1],
       \regs68H[6] [0]}), .in_7 ({\regs68H[7] [15], \regs68H[7] [14],
       \regs68H[7] [13], \regs68H[7] [12], \regs68H[7] [11],
       \regs68H[7] [10], \regs68H[7] [9], \regs68H[7] [8],
       \regs68H[7] [7], \regs68H[7] [6], \regs68H[7] [5],
       \regs68H[7] [4], \regs68H[7] [3], \regs68H[7] [2],
       \regs68H[7] [1], \regs68H[7] [0]}), .in_8 ({\regs68H[8] [15],
       \regs68H[8] [14], \regs68H[8] [13], \regs68H[8] [12],
       \regs68H[8] [11], \regs68H[8] [10], \regs68H[8] [9],
       \regs68H[8] [8], \regs68H[8] [7], \regs68H[8] [6],
       \regs68H[8] [5], \regs68H[8] [4], \regs68H[8] [3],
       \regs68H[8] [2], \regs68H[8] [1], \regs68H[8] [0]}), .in_9
       ({\regs68H[9] [15], \regs68H[9] [14], \regs68H[9] [13],
       \regs68H[9] [12], \regs68H[9] [11], \regs68H[9] [10],
       \regs68H[9] [9], \regs68H[9] [8], \regs68H[9] [7],
       \regs68H[9] [6], \regs68H[9] [5], \regs68H[9] [4],
       \regs68H[9] [3], \regs68H[9] [2], \regs68H[9] [1],
       \regs68H[9] [0]}), .in_10 ({\regs68H[10] [15], \regs68H[10]
       [14], \regs68H[10] [13], \regs68H[10] [12], \regs68H[10] [11],
       \regs68H[10] [10], \regs68H[10] [9], \regs68H[10] [8],
       \regs68H[10] [7], \regs68H[10] [6], \regs68H[10] [5],
       \regs68H[10] [4], \regs68H[10] [3], \regs68H[10] [2],
       \regs68H[10] [1], \regs68H[10] [0]}), .in_11 ({\regs68H[11]
       [15], \regs68H[11] [14], \regs68H[11] [13], \regs68H[11] [12],
       \regs68H[11] [11], \regs68H[11] [10], \regs68H[11] [9],
       \regs68H[11] [8], \regs68H[11] [7], \regs68H[11] [6],
       \regs68H[11] [5], \regs68H[11] [4], \regs68H[11] [3],
       \regs68H[11] [2], \regs68H[11] [1], \regs68H[11] [0]}), .in_12
       ({\regs68H[12] [15], \regs68H[12] [14], \regs68H[12] [13],
       \regs68H[12] [12], \regs68H[12] [11], \regs68H[12] [10],
       \regs68H[12] [9], \regs68H[12] [8], \regs68H[12] [7],
       \regs68H[12] [6], \regs68H[12] [5], \regs68H[12] [4],
       \regs68H[12] [3], \regs68H[12] [2], \regs68H[12] [1],
       \regs68H[12] [0]}), .in_13 ({\regs68H[13] [15], \regs68H[13]
       [14], \regs68H[13] [13], \regs68H[13] [12], \regs68H[13] [11],
       \regs68H[13] [10], \regs68H[13] [9], \regs68H[13] [8],
       \regs68H[13] [7], \regs68H[13] [6], \regs68H[13] [5],
       \regs68H[13] [4], \regs68H[13] [3], \regs68H[13] [2],
       \regs68H[13] [1], \regs68H[13] [0]}), .in_14 ({\regs68H[14]
       [15], \regs68H[14] [14], \regs68H[14] [13], \regs68H[14] [12],
       \regs68H[14] [11], \regs68H[14] [10], \regs68H[14] [9],
       \regs68H[14] [8], \regs68H[14] [7], \regs68H[14] [6],
       \regs68H[14] [5], \regs68H[14] [4], \regs68H[14] [3],
       \regs68H[14] [2], \regs68H[14] [1], \regs68H[14] [0]}), .in_15
       ({\regs68H[15] [15], \regs68H[15] [14], \regs68H[15] [13],
       \regs68H[15] [12], \regs68H[15] [11], \regs68H[15] [10],
       \regs68H[15] [9], \regs68H[15] [8], \regs68H[15] [7],
       \regs68H[15] [6], \regs68H[15] [5], \regs68H[15] [4],
       \regs68H[15] [3], \regs68H[15] [2], \regs68H[15] [1],
       \regs68H[15] [0]}), .in_16 ({\regs68H[16] [15], \regs68H[16]
       [14], \regs68H[16] [13], \regs68H[16] [12], \regs68H[16] [11],
       \regs68H[16] [10], \regs68H[16] [9], \regs68H[16] [8],
       \regs68H[16] [7], \regs68H[16] [6], \regs68H[16] [5],
       \regs68H[16] [4], \regs68H[16] [3], \regs68H[16] [2],
       \regs68H[16] [1], \regs68H[16] [0]}), .in_17 ({\regs68H[17]
       [15], \regs68H[17] [14], \regs68H[17] [13], \regs68H[17] [12],
       \regs68H[17] [11], \regs68H[17] [10], \regs68H[17] [9],
       \regs68H[17] [8], \regs68H[17] [7], \regs68H[17] [6],
       \regs68H[17] [5], \regs68H[17] [4], \regs68H[17] [3],
       \regs68H[17] [2], \regs68H[17] [1], \regs68H[17] [0]}), .z
       ({n_1075, n_1073, n_1071, n_1069, n_1067, n_1065, n_1063,
       n_1061, n_1059, n_1057, n_1055, n_1053, n_1051, n_1049, n_1047,
       n_1045}));
  fx68k_mux_2306 mux_abhMux_1357_10(.ctl ({Pch2Abh, \Nanod[rxh2abh] ,
       \Nanod[ryh2abh] , \Nanod[au2Ab] , \Nanod[aob2Ab] ,
       \Nanod[ath2Abh] }), .in_0 (PcH), .in_1 ({n_1074, n_1072, n_1070,
       n_1068, n_1066, n_1064, n_1062, n_1060, n_1058, n_1056, n_1054,
       n_1052, n_1050, n_1048, n_1046, n_1044}), .in_2 ({n_1075,
       n_1073, n_1071, n_1069, n_1067, n_1065, n_1063, n_1061, n_1059,
       n_1057, n_1055, n_1053, n_1051, n_1049, n_1047, n_1045}), .in_3
       (auReg[31:16]), .in_4 ({aob[31:24], eab[23:16]}), .in_5 (Ath),
       .z (abhMux));
  fx68k_bmux_1882 mux_1506_28(.ctl (\Nanod[dbl2rxl] ), .in_0 (AblOut),
       .in_1 (Dbl), .z ({n_1155, n_1153, n_1151, n_1149, n_1147,
       n_1145, n_1143, n_1141, n_1139, n_1137, n_1135, n_1133, n_1131,
       n_1129, n_1127, n_1125}));
  fx68k_bmux_1967 \mux_regs68L[actualRy]_1339_24 (.ctl (actualRy),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({n_1106, n_1104, n_1102, n_1100, n_1098, n_1096, n_1094,
       n_1092, n_1090, n_1088, n_1086, n_1084, n_1082, n_1080, n_1078,
       n_1076}));
  fx68k_bmux_1967 \mux_regs68L[actualRx]_1340_24 (.ctl (actualRx),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({n_1107, n_1105, n_1103, n_1101, n_1099, n_1097, n_1095,
       n_1093, n_1091, n_1089, n_1087, n_1085, n_1083, n_1081, n_1079,
       n_1077}));
  fx68k_mux_2324 mux_abdMux_1338_10(.ctl ({ryl2Abd, rxl2Abd,
       \Nanod[dbin2Abd] , \Nanod[alu2Abd] }), .in_0 ({n_1106, n_1104,
       n_1102, n_1100, n_1098, n_1096, n_1094, n_1092, n_1090, n_1088,
       n_1086, n_1084, n_1082, n_1080, n_1078, n_1076}), .in_1
       ({n_1107, n_1105, n_1103, n_1101, n_1099, n_1097, n_1095,
       n_1093, n_1091, n_1089, n_1087, n_1085, n_1083, n_1081, n_1079,
       n_1077}), .in_2 (dbin), .in_3 (aluOut), .z (abdMux));
  fx68k_bmux_1882 mux_1401_31(.ctl (ablIdle), .in_0 (preAbl), .in_1
       (preAbh), .z ({n_1123, n_1122, n_1121, n_1120, n_1119, n_1118,
       n_1117, n_1116, n_1115, n_1114, n_1113, n_1112, n_1111, n_1110,
       n_1109, n_1108}));
  fx68k_bmux_1882 mux_1401_11(.ctl (n_536), .in_0 ({n_1123, n_1122,
       n_1121, n_1120, n_1119, n_1118, n_1117, n_1116, n_1115, n_1114,
       n_1113, n_1112, n_1111, n_1110, n_1109, n_1108}), .in_1
       (preAbd), .z ({n_4258, n_4257, n_4256, n_4255, n_4254, n_4253,
       n_4252, n_4251, n_4250, n_4249, n_4248, n_4247, n_4246, n_4245,
       n_4244, n_4243}));
  fx68k_bmux_1882 \mux_regs68L[0]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_1154,
       n_1152, n_1150, n_1148, n_1146, n_1144, n_1142, n_1140, n_1138,
       n_1136, n_1134, n_1132, n_1130, n_1128, n_1126, n_1124}));
  fx68k_bmux_1882 \mux_regs68L[0]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_1154, n_1152, n_1150, n_1148, n_1146, n_1144, n_1142,
       n_1140, n_1138, n_1136, n_1134, n_1132, n_1130, n_1128, n_1126,
       n_1124}), .z ({n_1173, n_1172, n_1171, n_1170, n_1169, n_1168,
       n_1167, n_1166, n_1165, n_1164, n_1163, n_1162, n_1161, n_1160,
       n_1159, n_1158}));
  fx68k_mux_1995 \mux_regs68L[0]_1511_27 (.ctl ({n_669, n_670}), .in_0
       (Dbd), .in_1 ({n_1173, n_1172, n_1171, n_1170, n_1169, n_1168,
       n_1167, n_1166, n_1165, n_1164, n_1163, n_1162, n_1161, n_1160,
       n_1159, n_1158}), .z ({n_3999, n_3997, n_3995, n_3993, n_3991,
       n_3989, n_3987, n_3985, n_3983, n_3981, n_3979, n_3977, n_3975,
       n_3973, n_3971, n_3969}));
  fx68k_mux_1995 \mux_regs68L[0]_1513_16 (.ctl ({n_669, n_670}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_1173, n_1172, n_1171,
       n_1170, n_1169, n_1168, n_1167, n_1166, n_1165, n_1164, n_1163,
       n_1162, n_1161, n_1160, n_1159, n_1158}), .z ({n_3968, n_3967,
       n_3966, n_3965, n_3964, n_3963, n_3962, n_3961, n_3960, n_3958,
       n_3956, n_3954, n_3952, n_3950, n_3948, n_3946}));
  fx68k_bmux_1967 \mux_regs68L[actualRx]_1320_24 (.ctl (actualRx),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({n_1206, n_1204, n_1202, n_1200, n_1198, n_1196, n_1194,
       n_1192, n_1190, n_1188, n_1186, n_1184, n_1182, n_1180, n_1178,
       n_1176}));
  fx68k_bmux_1967 \mux_regs68L[actualRy]_1321_24 (.ctl (actualRy),
       .in_0 ({\regs68L[0] [15], \regs68L[0] [14], \regs68L[0] [13],
       \regs68L[0] [12], \regs68L[0] [11], \regs68L[0] [10],
       \regs68L[0] [9], \regs68L[0] [8], \regs68L[0] [7],
       \regs68L[0] [6], \regs68L[0] [5], \regs68L[0] [4],
       \regs68L[0] [3], \regs68L[0] [2], \regs68L[0] [1],
       \regs68L[0] [0]}), .in_1 ({\regs68L[1] [15], \regs68L[1] [14],
       \regs68L[1] [13], \regs68L[1] [12], \regs68L[1] [11],
       \regs68L[1] [10], \regs68L[1] [9], \regs68L[1] [8],
       \regs68L[1] [7], \regs68L[1] [6], \regs68L[1] [5],
       \regs68L[1] [4], \regs68L[1] [3], \regs68L[1] [2],
       \regs68L[1] [1], \regs68L[1] [0]}), .in_2 ({\regs68L[2] [15],
       \regs68L[2] [14], \regs68L[2] [13], \regs68L[2] [12],
       \regs68L[2] [11], \regs68L[2] [10], \regs68L[2] [9],
       \regs68L[2] [8], \regs68L[2] [7], \regs68L[2] [6],
       \regs68L[2] [5], \regs68L[2] [4], \regs68L[2] [3],
       \regs68L[2] [2], \regs68L[2] [1], \regs68L[2] [0]}), .in_3
       ({\regs68L[3] [15], \regs68L[3] [14], \regs68L[3] [13],
       \regs68L[3] [12], \regs68L[3] [11], \regs68L[3] [10],
       \regs68L[3] [9], \regs68L[3] [8], \regs68L[3] [7],
       \regs68L[3] [6], \regs68L[3] [5], \regs68L[3] [4],
       \regs68L[3] [3], \regs68L[3] [2], \regs68L[3] [1],
       \regs68L[3] [0]}), .in_4 ({\regs68L[4] [15], \regs68L[4] [14],
       \regs68L[4] [13], \regs68L[4] [12], \regs68L[4] [11],
       \regs68L[4] [10], \regs68L[4] [9], \regs68L[4] [8],
       \regs68L[4] [7], \regs68L[4] [6], \regs68L[4] [5],
       \regs68L[4] [4], \regs68L[4] [3], \regs68L[4] [2],
       \regs68L[4] [1], \regs68L[4] [0]}), .in_5 ({\regs68L[5] [15],
       \regs68L[5] [14], \regs68L[5] [13], \regs68L[5] [12],
       \regs68L[5] [11], \regs68L[5] [10], \regs68L[5] [9],
       \regs68L[5] [8], \regs68L[5] [7], \regs68L[5] [6],
       \regs68L[5] [5], \regs68L[5] [4], \regs68L[5] [3],
       \regs68L[5] [2], \regs68L[5] [1], \regs68L[5] [0]}), .in_6
       ({\regs68L[6] [15], \regs68L[6] [14], \regs68L[6] [13],
       \regs68L[6] [12], \regs68L[6] [11], \regs68L[6] [10],
       \regs68L[6] [9], \regs68L[6] [8], \regs68L[6] [7],
       \regs68L[6] [6], \regs68L[6] [5], \regs68L[6] [4],
       \regs68L[6] [3], \regs68L[6] [2], \regs68L[6] [1],
       \regs68L[6] [0]}), .in_7 ({\regs68L[7] [15], \regs68L[7] [14],
       \regs68L[7] [13], \regs68L[7] [12], \regs68L[7] [11],
       \regs68L[7] [10], \regs68L[7] [9], \regs68L[7] [8],
       \regs68L[7] [7], \regs68L[7] [6], \regs68L[7] [5],
       \regs68L[7] [4], \regs68L[7] [3], \regs68L[7] [2],
       \regs68L[7] [1], \regs68L[7] [0]}), .in_8 ({\regs68L[8] [15],
       \regs68L[8] [14], \regs68L[8] [13], \regs68L[8] [12],
       \regs68L[8] [11], \regs68L[8] [10], \regs68L[8] [9],
       \regs68L[8] [8], \regs68L[8] [7], \regs68L[8] [6],
       \regs68L[8] [5], \regs68L[8] [4], \regs68L[8] [3],
       \regs68L[8] [2], \regs68L[8] [1], \regs68L[8] [0]}), .in_9
       ({\regs68L[9] [15], \regs68L[9] [14], \regs68L[9] [13],
       \regs68L[9] [12], \regs68L[9] [11], \regs68L[9] [10],
       \regs68L[9] [9], \regs68L[9] [8], \regs68L[9] [7],
       \regs68L[9] [6], \regs68L[9] [5], \regs68L[9] [4],
       \regs68L[9] [3], \regs68L[9] [2], \regs68L[9] [1],
       \regs68L[9] [0]}), .in_10 ({\regs68L[10] [15], \regs68L[10]
       [14], \regs68L[10] [13], \regs68L[10] [12], \regs68L[10] [11],
       \regs68L[10] [10], \regs68L[10] [9], \regs68L[10] [8],
       \regs68L[10] [7], \regs68L[10] [6], \regs68L[10] [5],
       \regs68L[10] [4], \regs68L[10] [3], \regs68L[10] [2],
       \regs68L[10] [1], \regs68L[10] [0]}), .in_11 ({\regs68L[11]
       [15], \regs68L[11] [14], \regs68L[11] [13], \regs68L[11] [12],
       \regs68L[11] [11], \regs68L[11] [10], \regs68L[11] [9],
       \regs68L[11] [8], \regs68L[11] [7], \regs68L[11] [6],
       \regs68L[11] [5], \regs68L[11] [4], \regs68L[11] [3],
       \regs68L[11] [2], \regs68L[11] [1], \regs68L[11] [0]}), .in_12
       ({\regs68L[12] [15], \regs68L[12] [14], \regs68L[12] [13],
       \regs68L[12] [12], \regs68L[12] [11], \regs68L[12] [10],
       \regs68L[12] [9], \regs68L[12] [8], \regs68L[12] [7],
       \regs68L[12] [6], \regs68L[12] [5], \regs68L[12] [4],
       \regs68L[12] [3], \regs68L[12] [2], \regs68L[12] [1],
       \regs68L[12] [0]}), .in_13 ({\regs68L[13] [15], \regs68L[13]
       [14], \regs68L[13] [13], \regs68L[13] [12], \regs68L[13] [11],
       \regs68L[13] [10], \regs68L[13] [9], \regs68L[13] [8],
       \regs68L[13] [7], \regs68L[13] [6], \regs68L[13] [5],
       \regs68L[13] [4], \regs68L[13] [3], \regs68L[13] [2],
       \regs68L[13] [1], \regs68L[13] [0]}), .in_14 ({\regs68L[14]
       [15], \regs68L[14] [14], \regs68L[14] [13], \regs68L[14] [12],
       \regs68L[14] [11], \regs68L[14] [10], \regs68L[14] [9],
       \regs68L[14] [8], \regs68L[14] [7], \regs68L[14] [6],
       \regs68L[14] [5], \regs68L[14] [4], \regs68L[14] [3],
       \regs68L[14] [2], \regs68L[14] [1], \regs68L[14] [0]}), .in_15
       ({\regs68L[15] [15], \regs68L[15] [14], \regs68L[15] [13],
       \regs68L[15] [12], \regs68L[15] [11], \regs68L[15] [10],
       \regs68L[15] [9], \regs68L[15] [8], \regs68L[15] [7],
       \regs68L[15] [6], \regs68L[15] [5], \regs68L[15] [4],
       \regs68L[15] [3], \regs68L[15] [2], \regs68L[15] [1],
       \regs68L[15] [0]}), .in_16 ({\regs68L[16] [15], \regs68L[16]
       [14], \regs68L[16] [13], \regs68L[16] [12], \regs68L[16] [11],
       \regs68L[16] [10], \regs68L[16] [9], \regs68L[16] [8],
       \regs68L[16] [7], \regs68L[16] [6], \regs68L[16] [5],
       \regs68L[16] [4], \regs68L[16] [3], \regs68L[16] [2],
       \regs68L[16] [1], \regs68L[16] [0]}), .in_17 ({\regs68L[17]
       [15], \regs68L[17] [14], \regs68L[17] [13], \regs68L[17] [12],
       \regs68L[17] [11], \regs68L[17] [10], \regs68L[17] [9],
       \regs68L[17] [8], \regs68L[17] [7], \regs68L[17] [6],
       \regs68L[17] [5], \regs68L[17] [4], \regs68L[17] [3],
       \regs68L[17] [2], \regs68L[17] [1], \regs68L[17] [0]}), .z
       ({n_1207, n_1205, n_1203, n_1201, n_1199, n_1197, n_1195,
       n_1193, n_1191, n_1189, n_1187, n_1185, n_1183, n_1181, n_1179,
       n_1177}));
  fx68k_mux_2306 mux_dblMux_1319_10(.ctl ({rxl2Dbl, ryl2Dbl,
       \Nanod[ftu2Dbl] , \Nanod[au2Db] , \Nanod[atl2Dbl] , Pcl2Dbl}),
       .in_0 ({n_1206, n_1204, n_1202, n_1200, n_1198, n_1196, n_1194,
       n_1192, n_1190, n_1188, n_1186, n_1184, n_1182, n_1180, n_1178,
       n_1176}), .in_1 ({n_1207, n_1205, n_1203, n_1201, n_1199,
       n_1197, n_1195, n_1193, n_1191, n_1189, n_1187, n_1185, n_1183,
       n_1181, n_1179, n_1177}), .in_2 (ftu), .in_3 (auReg[15:0]),
       .in_4 (Atl), .in_5 (PcL), .z (dblMux));
  fx68k_bmux_1882 mux_1413_12(.ctl (\Nanod[dblDbh] ), .in_0 (preDbd),
       .in_1 (preDbh), .z ({n_1224, n_1223, n_1222, n_1221, n_1220,
       n_1219, n_1218, n_1217, n_1216, n_1215, n_1214, n_1213, n_1212,
       n_1211, n_1210, n_1209}));
  fx68k_bmux_1882 mux_Dbl_1410_8(.ctl (n_518), .in_0 ({n_1224, n_1223,
       n_1222, n_1221, n_1220, n_1219, n_1218, n_1217, n_1216, n_1215,
       n_1214, n_1213, n_1212, n_1211, n_1210, n_1209}), .in_1
       (preDbl), .z ({n_4210, n_4209, n_4208, n_4207, n_4206, n_4205,
       n_4204, n_4203, n_4202, n_4201, n_4200, n_4199, n_4198, n_4197,
       n_4196, n_4195}));
  fx68k_bmux_1520 mux_1462_38(.ctl (n_1226), .in_0 (2'b10), .in_1
       (2'b01), .z ({n_1233, n_1231}));
  fx68k_bmux_1503 mux_1468_38(.ctl (n_1226), .in_0 (1'b0), .in_1
       (1'b1), .z (n_1232));
  fx68k_bmux_2394 mux_auInpMux_1460_16(.ctl (\Nanod[auCntrl] ), .in_0
       (32'b00000000000000000000000000000000), .in_1
       ({30'b000000000000000000000000000000, n_1233, n_1231}), .in_2
       (32'b11111111111111111111111111111100), .in_3 ({Abh, AblOut}),
       .in_4 (32'b00000000000000000000000000000010), .in_5
       (32'b00000000000000000000000000000100), .in_6
       (32'b11111111111111111111111111111110), .in_7
       ({31'b1111111111111111111111111111111, n_1232}), .z (auInpMux));
  fx68k_bmux_1840 mux_auReg_1484_7(.ctl (\Clks[pwrUp] ), .in_0
       ({n_1265, n_1264, n_1263, n_1262, n_1261, n_1260, n_1259,
       n_1258, n_1257, n_1256, n_1255, n_1254, n_1253, n_1252, n_1251,
       n_1250, n_1249, n_1248, n_1247, n_1246, n_1245, n_1244, n_1243,
       n_1242, n_1241, n_1240, n_1239, n_1238, n_1237, n_1236, n_1235,
       n_1234}), .in_1 (32'b00000000000000000000000000000000), .z
       ({UNCONNECTED481, UNCONNECTED480, UNCONNECTED479,
       UNCONNECTED478, UNCONNECTED477, UNCONNECTED476, UNCONNECTED475,
       UNCONNECTED474, UNCONNECTED473, UNCONNECTED472, UNCONNECTED471,
       UNCONNECTED470, UNCONNECTED469, UNCONNECTED468, UNCONNECTED467,
       UNCONNECTED466, UNCONNECTED465, UNCONNECTED464, UNCONNECTED463,
       UNCONNECTED462, UNCONNECTED461, UNCONNECTED460, UNCONNECTED459,
       UNCONNECTED458, UNCONNECTED457, UNCONNECTED456, UNCONNECTED455,
       UNCONNECTED454, UNCONNECTED453, UNCONNECTED452, UNCONNECTED451,
       UNCONNECTED450}));
  fx68k_bmux_1882 mux_1443_22(.ctl (n_518), .in_0 (preDbd), .in_1
       (preDbl), .z ({n_1300, n_1298, n_1296, n_1294, n_1292, n_1290,
       n_1288, n_1286, n_1284, n_1282, n_1280, n_1278, n_1276, n_1274,
       n_1272, n_1270}));
  fx68k_bmux_1882 mux_1445_22(.ctl (n_552), .in_0 (preAbd), .in_1
       (preAbl), .z ({n_1301, n_1299, n_1297, n_1295, n_1293, n_1291,
       n_1289, n_1287, n_1285, n_1283, n_1281, n_1279, n_1277, n_1275,
       n_1273, n_1271}));
  fx68k_bmux_1840 mux_aob_1442_8(.ctl (\Nanod[db2Aob] ), .in_0
       ({preAbh, n_1301, n_1299, n_1297, n_1295, n_1293, n_1291,
       n_1289, n_1287, n_1285, n_1283, n_1281, n_1279, n_1277, n_1275,
       n_1273, n_1271}), .in_1 ({preDbh, n_1300, n_1298, n_1296,
       n_1294, n_1292, n_1290, n_1288, n_1286, n_1284, n_1282, n_1280,
       n_1278, n_1276, n_1274, n_1272, n_1270}), .z ({n_1333, n_1332,
       n_1331, n_1330, n_1329, n_1328, n_1327, n_1326, n_1325, n_1324,
       n_1323, n_1322, n_1321, n_1320, n_1319, n_1318, n_1317, n_1316,
       n_1315, n_1314, n_1313, n_1312, n_1311, n_1310, n_1309, n_1308,
       n_1307, n_1306, n_1305, n_1304, n_1303, n_1302}));
  fx68k_bmux_1840 mux_aob_1439_12(.ctl (n_451), .in_0 ({n_1333, n_1332,
       n_1331, n_1330, n_1329, n_1328, n_1327, n_1326, n_1325, n_1324,
       n_1323, n_1322, n_1321, n_1320, n_1319, n_1318, n_1317, n_1316,
       n_1315, n_1314, n_1313, n_1312, n_1311, n_1310, n_1309, n_1308,
       n_1307, n_1306, n_1305, n_1304, n_1303, n_1302}), .in_1 (auReg),
       .z ({n_4314, n_4313, n_4312, n_4311, n_4310, n_4309, n_4308,
       n_4307, n_4306, n_4305, n_4304, n_4303, n_4302, n_4301, n_4300,
       n_4299, n_4298, n_4297, n_4296, n_4295, n_4294, n_4293, n_4292,
       n_4291, n_4290, n_4289, n_4288, n_4287, n_4286, n_4285, n_4284,
       n_4282}));
  fx68k_bmux_1883 mux_dobInput_1647_16(.ctl (\Nanod[dobCtrl] ), .in_0
       ({_X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_, _X_,
       _X_, _X_, _X_, _X_}), .in_1 (Dbd), .in_2 ({Abd[15:3],
       dcrInput[2:0]}), .in_3 (aluOut), .z (dobInput));
  fx68k_bmux_1504 mux_1263_12(.ctl (\Nanod[rz] ), .in_0
       ({\Irdecod[ryIsAreg] , \Irdecod[ry] }), .in_1 (Irc[15:12]), .z
       (ryReg));
  fx68k_bmux_1503 mux_ryIsSp_1257_22(.ctl (n_449), .in_0 (n_1344),
       .in_1 (1'b0), .z (ryIsSp));
  fx68k_mux_1959 mux_dbdIdle_1309_10(.ctl ({ryl2Dbd, rxl2Dbd,
       \Nanod[alue2Dbd] , \Nanod[dbin2Dbd] , \Nanod[alu2Dbd] ,
       \Nanod[dcr2Dbd] , n_1357}), .in_0 (1'b0), .in_1 (1'b0), .in_2
       (1'b0), .in_3 (1'b0), .in_4 (1'b0), .in_5 (1'b0), .in_6 (1'b1),
       .z (dbdIdle));
  fx68k_bmux_1882 mux_1415_30(.ctl (dblIdle), .in_0 (preDbl), .in_1
       (preDbh), .z ({n_1374, n_1373, n_1372, n_1371, n_1370, n_1369,
       n_1368, n_1367, n_1366, n_1365, n_1364, n_1363, n_1362, n_1361,
       n_1360, n_1359}));
  fx68k_bmux_1882 mux_1415_11(.ctl (n_1358), .in_0 ({n_1374, n_1373,
       n_1372, n_1371, n_1370, n_1369, n_1368, n_1367, n_1366, n_1365,
       n_1364, n_1363, n_1362, n_1361, n_1360, n_1359}), .in_1
       (preDbd), .z ({n_4274, n_4273, n_4272, n_4271, n_4270, n_4269,
       n_4268, n_4267, n_4266, n_4265, n_4264, n_4263, n_4262, n_4261,
       n_4260, n_4259}));
  fx68k_bmux_1882 mux_alub_1632_8(.ctl (\Nanod[dbd2Alub] ), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_6307, n_6306,
       n_6305, n_6304, n_6303, n_6302, n_6301, n_6300, n_6299, n_6298,
       n_6297, n_6296, n_6295, n_6294, n_6293, n_6291}));
  fx68k_bmux_1503 mux_dcr4_1618_7(.ctl (\Clks[pwrUp] ), .in_0 (Abd[4]),
       .in_1 (1'b0), .z (UNCONNECTED482));
  fx68k_bmux_1854 mux_ryMux_1265_15(.ctl (n_523), .in_0 ({1'b0,
       ryReg}), .in_1 (5'b10000), .z ({n_1380, n_1379, n_1378, n_1377,
       n_1376}));
  fx68k_bmux_1854 mux_ryMux_1257_22(.ctl (n_449), .in_0 ({n_1380,
       n_1379, n_1378, n_1377, n_1376}), .in_1 (5'b10001), .z (ryMux));
  fx68k_bmux_1882 \mux_regs68L[1]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_3814,
       n_3813, n_3812, n_3811, n_3810, n_3809, n_3808, n_3807, n_3806,
       n_3805, n_3804, n_3803, n_3802, n_3801, n_3800, n_3799}));
  fx68k_bmux_1882 \mux_regs68L[2]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_1396,
       n_1395, n_1394, n_1393, n_1392, n_1391, n_1390, n_1389, n_1388,
       n_1387, n_1386, n_1385, n_1384, n_1383, n_1382, n_1381}));
  fx68k_bmux_1882 \mux_regs68L[2]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_1396, n_1395, n_1394, n_1393, n_1392, n_1391, n_1390,
       n_1389, n_1388, n_1387, n_1386, n_1385, n_1384, n_1383, n_1382,
       n_1381}), .z ({n_1414, n_1413, n_1412, n_1411, n_1410, n_1409,
       n_1408, n_1407, n_1406, n_1405, n_1404, n_1403, n_1402, n_1401,
       n_1400, n_1399}));
  fx68k_mux_1995 \mux_regs68L[2]_1511_27 (.ctl ({n_737, n_738}), .in_0
       (Dbd), .in_1 ({n_1414, n_1413, n_1412, n_1411, n_1410, n_1409,
       n_1408, n_1407, n_1406, n_1405, n_1404, n_1403, n_1402, n_1401,
       n_1400, n_1399}), .z ({n_1473, n_1471, n_1469, n_1467, n_1465,
       n_1463, n_1461, n_1459, n_1457, n_1455, n_1453, n_1451, n_1449,
       n_1447, n_1445, n_1443}));
  fx68k_mux_2428 \mux_regs68L[2]_1512_28 (.ctl ({n_737, n_738}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_1406, n_1405, n_1404,
       n_1403, n_1402, n_1401, n_1400, n_1399}), .z ({n_1433, n_1431,
       n_1429, n_1427, n_1425, n_1423, n_1421, n_1419}));
  fx68k_mux_1995 \mux_regs68L[2]_1513_16 (.ctl ({n_737, n_738}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_1414, n_1413, n_1412,
       n_1411, n_1410, n_1409, n_1408, n_1407, n_1406, n_1405, n_1404,
       n_1403, n_1402, n_1401, n_1400, n_1399}), .z ({n_1442, n_1441,
       n_1440, n_1439, n_1438, n_1437, n_1436, n_1435, n_1434, n_1432,
       n_1430, n_1428, n_1426, n_1424, n_1422, n_1420}));
  fx68k_bmux_1882 \mux_regs68L[2]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_1442, n_1441, n_1440, n_1439, n_1438, n_1437, n_1436,
       n_1435, n_1434, n_1432, n_1430, n_1428, n_1426, n_1424, n_1422,
       n_1420}), .in_1 ({n_1414, n_1413, n_1412, n_1411, n_1410,
       n_1409, n_1408, n_1407, n_1433, n_1431, n_1429, n_1427, n_1425,
       n_1423, n_1421, n_1419}), .z ({n_1474, n_1472, n_1470, n_1468,
       n_1466, n_1464, n_1462, n_1460, n_1458, n_1456, n_1454, n_1452,
       n_1450, n_1448, n_1446, n_1444}));
  fx68k_bmux_1882 \mux_regs68L[2]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_1474, n_1472, n_1470, n_1468, n_1466, n_1464, n_1462,
       n_1460, n_1458, n_1456, n_1454, n_1452, n_1450, n_1448, n_1446,
       n_1444}), .in_1 ({n_1473, n_1471, n_1469, n_1467, n_1465,
       n_1463, n_1461, n_1459, n_1457, n_1455, n_1453, n_1451, n_1449,
       n_1447, n_1445, n_1443}), .z ({n_1523, n_1521, n_1519, n_1517,
       n_1515, n_1513, n_1511, n_1509, n_1507, n_1505, n_1503, n_1501,
       n_1499, n_1497, n_1495, n_1493}));
  fx68k_bmux_1882 mux_1516_28(.ctl (\Nanod[dbl2ryl] ), .in_0 (AblOut),
       .in_1 (Dbl), .z ({n_1492, n_1491, n_1490, n_1489, n_1488,
       n_1487, n_1486, n_1485, n_1484, n_1483, n_1482, n_1481, n_1480,
       n_1479, n_1478, n_1477}));
  fx68k_mux_1995 \mux_regs68L[2]_1516_6 (.ctl ({n_737, n_738}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_1414, n_1413, n_1412, n_1411, n_1410,
       n_1409, n_1408, n_1407, n_1406, n_1405, n_1404, n_1403, n_1402,
       n_1401, n_1400, n_1399}), .z ({n_1524, n_1522, n_1520, n_1518,
       n_1516, n_1514, n_1512, n_1510, n_1508, n_1506, n_1504, n_1502,
       n_1500, n_1498, n_1496, n_1494}));
  fx68k_bmux_1882 \mux_regs68L[2]_1510_9 (.ctl (n_521), .in_0 ({n_1524,
       n_1522, n_1520, n_1518, n_1516, n_1514, n_1512, n_1510, n_1508,
       n_1506, n_1504, n_1502, n_1500, n_1498, n_1496, n_1494}), .in_1
       ({n_1523, n_1521, n_1519, n_1517, n_1515, n_1513, n_1511,
       n_1509, n_1507, n_1505, n_1503, n_1501, n_1499, n_1497, n_1495,
       n_1493}), .z ({n_1540, n_1539, n_1538, n_1537, n_1536, n_1535,
       n_1534, n_1533, n_1532, n_1531, n_1530, n_1529, n_1528, n_1527,
       n_1526, n_1525}));
  fx68k_bmux_1882 \mux_regs68L[2]_1509_22 (.ctl (n_520), .in_0
       ({n_1414, n_1413, n_1412, n_1411, n_1410, n_1409, n_1408,
       n_1407, n_1406, n_1405, n_1404, n_1403, n_1402, n_1401, n_1400,
       n_1399}), .in_1 ({n_1540, n_1539, n_1538, n_1537, n_1536,
       n_1535, n_1534, n_1533, n_1532, n_1531, n_1530, n_1529, n_1528,
       n_1527, n_1526, n_1525}), .z ({n_5584, n_5583, n_5582, n_5581,
       n_5580, n_5579, n_5578, n_5576, n_5575, n_5574, n_5573, n_5572,
       n_5571, n_5570, n_5569, n_5567}));
  fx68k_bmux_1882 \mux_regs68L[3]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_1556,
       n_1555, n_1554, n_1553, n_1552, n_1551, n_1550, n_1549, n_1548,
       n_1547, n_1546, n_1545, n_1544, n_1543, n_1542, n_1541}));
  fx68k_bmux_1882 \mux_regs68L[3]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_1556, n_1555, n_1554, n_1553, n_1552, n_1551, n_1550,
       n_1549, n_1548, n_1547, n_1546, n_1545, n_1544, n_1543, n_1542,
       n_1541}), .z ({n_1574, n_1573, n_1572, n_1571, n_1570, n_1569,
       n_1568, n_1567, n_1566, n_1565, n_1564, n_1563, n_1562, n_1561,
       n_1560, n_1559}));
  fx68k_mux_1995 \mux_regs68L[3]_1511_27 (.ctl ({n_755, n_756}), .in_0
       (Dbd), .in_1 ({n_1574, n_1573, n_1572, n_1571, n_1570, n_1569,
       n_1568, n_1567, n_1566, n_1565, n_1564, n_1563, n_1562, n_1561,
       n_1560, n_1559}), .z ({n_1633, n_1631, n_1629, n_1627, n_1625,
       n_1623, n_1621, n_1619, n_1617, n_1615, n_1613, n_1611, n_1609,
       n_1607, n_1605, n_1603}));
  fx68k_mux_2428 \mux_regs68L[3]_1512_28 (.ctl ({n_755, n_756}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_1566, n_1565, n_1564,
       n_1563, n_1562, n_1561, n_1560, n_1559}), .z ({n_1593, n_1591,
       n_1589, n_1587, n_1585, n_1583, n_1581, n_1579}));
  fx68k_mux_1995 \mux_regs68L[3]_1513_16 (.ctl ({n_755, n_756}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_1574, n_1573, n_1572,
       n_1571, n_1570, n_1569, n_1568, n_1567, n_1566, n_1565, n_1564,
       n_1563, n_1562, n_1561, n_1560, n_1559}), .z ({n_1602, n_1601,
       n_1600, n_1599, n_1598, n_1597, n_1596, n_1595, n_1594, n_1592,
       n_1590, n_1588, n_1586, n_1584, n_1582, n_1580}));
  fx68k_bmux_1882 \mux_regs68L[3]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_1602, n_1601, n_1600, n_1599, n_1598, n_1597, n_1596,
       n_1595, n_1594, n_1592, n_1590, n_1588, n_1586, n_1584, n_1582,
       n_1580}), .in_1 ({n_1574, n_1573, n_1572, n_1571, n_1570,
       n_1569, n_1568, n_1567, n_1593, n_1591, n_1589, n_1587, n_1585,
       n_1583, n_1581, n_1579}), .z ({n_1634, n_1632, n_1630, n_1628,
       n_1626, n_1624, n_1622, n_1620, n_1618, n_1616, n_1614, n_1612,
       n_1610, n_1608, n_1606, n_1604}));
  fx68k_bmux_1882 \mux_regs68L[3]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_1634, n_1632, n_1630, n_1628, n_1626, n_1624, n_1622,
       n_1620, n_1618, n_1616, n_1614, n_1612, n_1610, n_1608, n_1606,
       n_1604}), .in_1 ({n_1633, n_1631, n_1629, n_1627, n_1625,
       n_1623, n_1621, n_1619, n_1617, n_1615, n_1613, n_1611, n_1609,
       n_1607, n_1605, n_1603}), .z ({n_1667, n_1665, n_1663, n_1661,
       n_1659, n_1657, n_1655, n_1653, n_1651, n_1649, n_1647, n_1645,
       n_1643, n_1641, n_1639, n_1637}));
  fx68k_mux_1995 \mux_regs68L[3]_1516_6 (.ctl ({n_755, n_756}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_1574, n_1573, n_1572, n_1571, n_1570,
       n_1569, n_1568, n_1567, n_1566, n_1565, n_1564, n_1563, n_1562,
       n_1561, n_1560, n_1559}), .z ({n_1668, n_1666, n_1664, n_1662,
       n_1660, n_1658, n_1656, n_1654, n_1652, n_1650, n_1648, n_1646,
       n_1644, n_1642, n_1640, n_1638}));
  fx68k_bmux_1882 \mux_regs68L[3]_1510_9 (.ctl (n_521), .in_0 ({n_1668,
       n_1666, n_1664, n_1662, n_1660, n_1658, n_1656, n_1654, n_1652,
       n_1650, n_1648, n_1646, n_1644, n_1642, n_1640, n_1638}), .in_1
       ({n_1667, n_1665, n_1663, n_1661, n_1659, n_1657, n_1655,
       n_1653, n_1651, n_1649, n_1647, n_1645, n_1643, n_1641, n_1639,
       n_1637}), .z ({n_1684, n_1683, n_1682, n_1681, n_1680, n_1679,
       n_1678, n_1677, n_1676, n_1675, n_1674, n_1673, n_1672, n_1671,
       n_1670, n_1669}));
  fx68k_bmux_1882 \mux_regs68L[3]_1509_22 (.ctl (n_520), .in_0
       ({n_1574, n_1573, n_1572, n_1571, n_1570, n_1569, n_1568,
       n_1567, n_1566, n_1565, n_1564, n_1563, n_1562, n_1561, n_1560,
       n_1559}), .in_1 ({n_1684, n_1683, n_1682, n_1681, n_1680,
       n_1679, n_1678, n_1677, n_1676, n_1675, n_1674, n_1673, n_1672,
       n_1671, n_1670, n_1669}), .z ({n_5505, n_5504, n_5503, n_5502,
       n_5501, n_5500, n_5499, n_5497, n_5496, n_5495, n_5494, n_5493,
       n_5492, n_5491, n_5490, n_5488}));
  fx68k_bmux_1882 \mux_regs68L[4]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_1700,
       n_1699, n_1698, n_1697, n_1696, n_1695, n_1694, n_1693, n_1692,
       n_1691, n_1690, n_1689, n_1688, n_1687, n_1686, n_1685}));
  fx68k_bmux_1882 \mux_regs68L[4]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_1700, n_1699, n_1698, n_1697, n_1696, n_1695, n_1694,
       n_1693, n_1692, n_1691, n_1690, n_1689, n_1688, n_1687, n_1686,
       n_1685}), .z ({n_1718, n_1717, n_1716, n_1715, n_1714, n_1713,
       n_1712, n_1711, n_1710, n_1709, n_1708, n_1707, n_1706, n_1705,
       n_1704, n_1703}));
  fx68k_mux_1995 \mux_regs68L[4]_1511_27 (.ctl ({n_773, n_774}), .in_0
       (Dbd), .in_1 ({n_1718, n_1717, n_1716, n_1715, n_1714, n_1713,
       n_1712, n_1711, n_1710, n_1709, n_1708, n_1707, n_1706, n_1705,
       n_1704, n_1703}), .z ({n_1777, n_1775, n_1773, n_1771, n_1769,
       n_1767, n_1765, n_1763, n_1761, n_1759, n_1757, n_1755, n_1753,
       n_1751, n_1749, n_1747}));
  fx68k_mux_2428 \mux_regs68L[4]_1512_28 (.ctl ({n_773, n_774}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_1710, n_1709, n_1708,
       n_1707, n_1706, n_1705, n_1704, n_1703}), .z ({n_1737, n_1735,
       n_1733, n_1731, n_1729, n_1727, n_1725, n_1723}));
  fx68k_mux_1995 \mux_regs68L[4]_1513_16 (.ctl ({n_773, n_774}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_1718, n_1717, n_1716,
       n_1715, n_1714, n_1713, n_1712, n_1711, n_1710, n_1709, n_1708,
       n_1707, n_1706, n_1705, n_1704, n_1703}), .z ({n_1746, n_1745,
       n_1744, n_1743, n_1742, n_1741, n_1740, n_1739, n_1738, n_1736,
       n_1734, n_1732, n_1730, n_1728, n_1726, n_1724}));
  fx68k_bmux_1882 \mux_regs68L[4]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_1746, n_1745, n_1744, n_1743, n_1742, n_1741, n_1740,
       n_1739, n_1738, n_1736, n_1734, n_1732, n_1730, n_1728, n_1726,
       n_1724}), .in_1 ({n_1718, n_1717, n_1716, n_1715, n_1714,
       n_1713, n_1712, n_1711, n_1737, n_1735, n_1733, n_1731, n_1729,
       n_1727, n_1725, n_1723}), .z ({n_1778, n_1776, n_1774, n_1772,
       n_1770, n_1768, n_1766, n_1764, n_1762, n_1760, n_1758, n_1756,
       n_1754, n_1752, n_1750, n_1748}));
  fx68k_bmux_1882 \mux_regs68L[4]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_1778, n_1776, n_1774, n_1772, n_1770, n_1768, n_1766,
       n_1764, n_1762, n_1760, n_1758, n_1756, n_1754, n_1752, n_1750,
       n_1748}), .in_1 ({n_1777, n_1775, n_1773, n_1771, n_1769,
       n_1767, n_1765, n_1763, n_1761, n_1759, n_1757, n_1755, n_1753,
       n_1751, n_1749, n_1747}), .z ({n_1811, n_1809, n_1807, n_1805,
       n_1803, n_1801, n_1799, n_1797, n_1795, n_1793, n_1791, n_1789,
       n_1787, n_1785, n_1783, n_1781}));
  fx68k_mux_1995 \mux_regs68L[4]_1516_6 (.ctl ({n_773, n_774}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_1718, n_1717, n_1716, n_1715, n_1714,
       n_1713, n_1712, n_1711, n_1710, n_1709, n_1708, n_1707, n_1706,
       n_1705, n_1704, n_1703}), .z ({n_1812, n_1810, n_1808, n_1806,
       n_1804, n_1802, n_1800, n_1798, n_1796, n_1794, n_1792, n_1790,
       n_1788, n_1786, n_1784, n_1782}));
  fx68k_bmux_1882 \mux_regs68L[4]_1510_9 (.ctl (n_521), .in_0 ({n_1812,
       n_1810, n_1808, n_1806, n_1804, n_1802, n_1800, n_1798, n_1796,
       n_1794, n_1792, n_1790, n_1788, n_1786, n_1784, n_1782}), .in_1
       ({n_1811, n_1809, n_1807, n_1805, n_1803, n_1801, n_1799,
       n_1797, n_1795, n_1793, n_1791, n_1789, n_1787, n_1785, n_1783,
       n_1781}), .z ({n_1828, n_1827, n_1826, n_1825, n_1824, n_1823,
       n_1822, n_1821, n_1820, n_1819, n_1818, n_1817, n_1816, n_1815,
       n_1814, n_1813}));
  fx68k_bmux_1882 \mux_regs68L[4]_1509_22 (.ctl (n_520), .in_0
       ({n_1718, n_1717, n_1716, n_1715, n_1714, n_1713, n_1712,
       n_1711, n_1710, n_1709, n_1708, n_1707, n_1706, n_1705, n_1704,
       n_1703}), .in_1 ({n_1828, n_1827, n_1826, n_1825, n_1824,
       n_1823, n_1822, n_1821, n_1820, n_1819, n_1818, n_1817, n_1816,
       n_1815, n_1814, n_1813}), .z ({n_5426, n_5425, n_5424, n_5423,
       n_5422, n_5421, n_5420, n_5418, n_5417, n_5416, n_5415, n_5414,
       n_5413, n_5412, n_5411, n_5409}));
  fx68k_bmux_1882 \mux_regs68L[5]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_1844,
       n_1843, n_1842, n_1841, n_1840, n_1839, n_1838, n_1837, n_1836,
       n_1835, n_1834, n_1833, n_1832, n_1831, n_1830, n_1829}));
  fx68k_bmux_1882 \mux_regs68L[5]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_1844, n_1843, n_1842, n_1841, n_1840, n_1839, n_1838,
       n_1837, n_1836, n_1835, n_1834, n_1833, n_1832, n_1831, n_1830,
       n_1829}), .z ({n_1862, n_1861, n_1860, n_1859, n_1858, n_1857,
       n_1856, n_1855, n_1854, n_1853, n_1852, n_1851, n_1850, n_1849,
       n_1848, n_1847}));
  fx68k_mux_1995 \mux_regs68L[5]_1511_27 (.ctl ({n_791, n_792}), .in_0
       (Dbd), .in_1 ({n_1862, n_1861, n_1860, n_1859, n_1858, n_1857,
       n_1856, n_1855, n_1854, n_1853, n_1852, n_1851, n_1850, n_1849,
       n_1848, n_1847}), .z ({n_1921, n_1919, n_1917, n_1915, n_1913,
       n_1911, n_1909, n_1907, n_1905, n_1903, n_1901, n_1899, n_1897,
       n_1895, n_1893, n_1891}));
  fx68k_mux_2428 \mux_regs68L[5]_1512_28 (.ctl ({n_791, n_792}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_1854, n_1853, n_1852,
       n_1851, n_1850, n_1849, n_1848, n_1847}), .z ({n_1881, n_1879,
       n_1877, n_1875, n_1873, n_1871, n_1869, n_1867}));
  fx68k_mux_1995 \mux_regs68L[5]_1513_16 (.ctl ({n_791, n_792}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_1862, n_1861, n_1860,
       n_1859, n_1858, n_1857, n_1856, n_1855, n_1854, n_1853, n_1852,
       n_1851, n_1850, n_1849, n_1848, n_1847}), .z ({n_1890, n_1889,
       n_1888, n_1887, n_1886, n_1885, n_1884, n_1883, n_1882, n_1880,
       n_1878, n_1876, n_1874, n_1872, n_1870, n_1868}));
  fx68k_bmux_1882 \mux_regs68L[5]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_1890, n_1889, n_1888, n_1887, n_1886, n_1885, n_1884,
       n_1883, n_1882, n_1880, n_1878, n_1876, n_1874, n_1872, n_1870,
       n_1868}), .in_1 ({n_1862, n_1861, n_1860, n_1859, n_1858,
       n_1857, n_1856, n_1855, n_1881, n_1879, n_1877, n_1875, n_1873,
       n_1871, n_1869, n_1867}), .z ({n_1922, n_1920, n_1918, n_1916,
       n_1914, n_1912, n_1910, n_1908, n_1906, n_1904, n_1902, n_1900,
       n_1898, n_1896, n_1894, n_1892}));
  fx68k_bmux_1882 \mux_regs68L[5]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_1922, n_1920, n_1918, n_1916, n_1914, n_1912, n_1910,
       n_1908, n_1906, n_1904, n_1902, n_1900, n_1898, n_1896, n_1894,
       n_1892}), .in_1 ({n_1921, n_1919, n_1917, n_1915, n_1913,
       n_1911, n_1909, n_1907, n_1905, n_1903, n_1901, n_1899, n_1897,
       n_1895, n_1893, n_1891}), .z ({n_1955, n_1953, n_1951, n_1949,
       n_1947, n_1945, n_1943, n_1941, n_1939, n_1937, n_1935, n_1933,
       n_1931, n_1929, n_1927, n_1925}));
  fx68k_mux_1995 \mux_regs68L[5]_1516_6 (.ctl ({n_791, n_792}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_1862, n_1861, n_1860, n_1859, n_1858,
       n_1857, n_1856, n_1855, n_1854, n_1853, n_1852, n_1851, n_1850,
       n_1849, n_1848, n_1847}), .z ({n_1956, n_1954, n_1952, n_1950,
       n_1948, n_1946, n_1944, n_1942, n_1940, n_1938, n_1936, n_1934,
       n_1932, n_1930, n_1928, n_1926}));
  fx68k_bmux_1882 \mux_regs68L[5]_1510_9 (.ctl (n_521), .in_0 ({n_1956,
       n_1954, n_1952, n_1950, n_1948, n_1946, n_1944, n_1942, n_1940,
       n_1938, n_1936, n_1934, n_1932, n_1930, n_1928, n_1926}), .in_1
       ({n_1955, n_1953, n_1951, n_1949, n_1947, n_1945, n_1943,
       n_1941, n_1939, n_1937, n_1935, n_1933, n_1931, n_1929, n_1927,
       n_1925}), .z ({n_1972, n_1971, n_1970, n_1969, n_1968, n_1967,
       n_1966, n_1965, n_1964, n_1963, n_1962, n_1961, n_1960, n_1959,
       n_1958, n_1957}));
  fx68k_bmux_1882 \mux_regs68L[5]_1509_22 (.ctl (n_520), .in_0
       ({n_1862, n_1861, n_1860, n_1859, n_1858, n_1857, n_1856,
       n_1855, n_1854, n_1853, n_1852, n_1851, n_1850, n_1849, n_1848,
       n_1847}), .in_1 ({n_1972, n_1971, n_1970, n_1969, n_1968,
       n_1967, n_1966, n_1965, n_1964, n_1963, n_1962, n_1961, n_1960,
       n_1959, n_1958, n_1957}), .z ({n_5347, n_5346, n_5345, n_5344,
       n_5343, n_5342, n_5341, n_5339, n_5338, n_5337, n_5336, n_5335,
       n_5334, n_5333, n_5332, n_5330}));
  fx68k_bmux_1882 \mux_regs68L[6]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_1988,
       n_1987, n_1986, n_1985, n_1984, n_1983, n_1982, n_1981, n_1980,
       n_1979, n_1978, n_1977, n_1976, n_1975, n_1974, n_1973}));
  fx68k_bmux_1882 \mux_regs68L[6]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_1988, n_1987, n_1986, n_1985, n_1984, n_1983, n_1982,
       n_1981, n_1980, n_1979, n_1978, n_1977, n_1976, n_1975, n_1974,
       n_1973}), .z ({n_2006, n_2005, n_2004, n_2003, n_2002, n_2001,
       n_2000, n_1999, n_1998, n_1997, n_1996, n_1995, n_1994, n_1993,
       n_1992, n_1991}));
  fx68k_mux_1995 \mux_regs68L[6]_1511_27 (.ctl ({n_809, n_810}), .in_0
       (Dbd), .in_1 ({n_2006, n_2005, n_2004, n_2003, n_2002, n_2001,
       n_2000, n_1999, n_1998, n_1997, n_1996, n_1995, n_1994, n_1993,
       n_1992, n_1991}), .z ({n_2065, n_2063, n_2061, n_2059, n_2057,
       n_2055, n_2053, n_2051, n_2049, n_2047, n_2045, n_2043, n_2041,
       n_2039, n_2037, n_2035}));
  fx68k_mux_2428 \mux_regs68L[6]_1512_28 (.ctl ({n_809, n_810}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_1998, n_1997, n_1996,
       n_1995, n_1994, n_1993, n_1992, n_1991}), .z ({n_2025, n_2023,
       n_2021, n_2019, n_2017, n_2015, n_2013, n_2011}));
  fx68k_mux_1995 \mux_regs68L[6]_1513_16 (.ctl ({n_809, n_810}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_2006, n_2005, n_2004,
       n_2003, n_2002, n_2001, n_2000, n_1999, n_1998, n_1997, n_1996,
       n_1995, n_1994, n_1993, n_1992, n_1991}), .z ({n_2034, n_2033,
       n_2032, n_2031, n_2030, n_2029, n_2028, n_2027, n_2026, n_2024,
       n_2022, n_2020, n_2018, n_2016, n_2014, n_2012}));
  fx68k_bmux_1882 \mux_regs68L[6]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_2034, n_2033, n_2032, n_2031, n_2030, n_2029, n_2028,
       n_2027, n_2026, n_2024, n_2022, n_2020, n_2018, n_2016, n_2014,
       n_2012}), .in_1 ({n_2006, n_2005, n_2004, n_2003, n_2002,
       n_2001, n_2000, n_1999, n_2025, n_2023, n_2021, n_2019, n_2017,
       n_2015, n_2013, n_2011}), .z ({n_2066, n_2064, n_2062, n_2060,
       n_2058, n_2056, n_2054, n_2052, n_2050, n_2048, n_2046, n_2044,
       n_2042, n_2040, n_2038, n_2036}));
  fx68k_bmux_1882 \mux_regs68L[6]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_2066, n_2064, n_2062, n_2060, n_2058, n_2056, n_2054,
       n_2052, n_2050, n_2048, n_2046, n_2044, n_2042, n_2040, n_2038,
       n_2036}), .in_1 ({n_2065, n_2063, n_2061, n_2059, n_2057,
       n_2055, n_2053, n_2051, n_2049, n_2047, n_2045, n_2043, n_2041,
       n_2039, n_2037, n_2035}), .z ({n_2099, n_2097, n_2095, n_2093,
       n_2091, n_2089, n_2087, n_2085, n_2083, n_2081, n_2079, n_2077,
       n_2075, n_2073, n_2071, n_2069}));
  fx68k_mux_1995 \mux_regs68L[6]_1516_6 (.ctl ({n_809, n_810}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_2006, n_2005, n_2004, n_2003, n_2002,
       n_2001, n_2000, n_1999, n_1998, n_1997, n_1996, n_1995, n_1994,
       n_1993, n_1992, n_1991}), .z ({n_2100, n_2098, n_2096, n_2094,
       n_2092, n_2090, n_2088, n_2086, n_2084, n_2082, n_2080, n_2078,
       n_2076, n_2074, n_2072, n_2070}));
  fx68k_bmux_1882 \mux_regs68L[6]_1510_9 (.ctl (n_521), .in_0 ({n_2100,
       n_2098, n_2096, n_2094, n_2092, n_2090, n_2088, n_2086, n_2084,
       n_2082, n_2080, n_2078, n_2076, n_2074, n_2072, n_2070}), .in_1
       ({n_2099, n_2097, n_2095, n_2093, n_2091, n_2089, n_2087,
       n_2085, n_2083, n_2081, n_2079, n_2077, n_2075, n_2073, n_2071,
       n_2069}), .z ({n_2116, n_2115, n_2114, n_2113, n_2112, n_2111,
       n_2110, n_2109, n_2108, n_2107, n_2106, n_2105, n_2104, n_2103,
       n_2102, n_2101}));
  fx68k_bmux_1882 \mux_regs68L[6]_1509_22 (.ctl (n_520), .in_0
       ({n_2006, n_2005, n_2004, n_2003, n_2002, n_2001, n_2000,
       n_1999, n_1998, n_1997, n_1996, n_1995, n_1994, n_1993, n_1992,
       n_1991}), .in_1 ({n_2116, n_2115, n_2114, n_2113, n_2112,
       n_2111, n_2110, n_2109, n_2108, n_2107, n_2106, n_2105, n_2104,
       n_2103, n_2102, n_2101}), .z ({n_5268, n_5267, n_5266, n_5265,
       n_5264, n_5263, n_5262, n_5260, n_5259, n_5258, n_5257, n_5256,
       n_5255, n_5254, n_5253, n_5251}));
  fx68k_bmux_1882 \mux_regs68L[7]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_2132,
       n_2131, n_2130, n_2129, n_2128, n_2127, n_2126, n_2125, n_2124,
       n_2123, n_2122, n_2121, n_2120, n_2119, n_2118, n_2117}));
  fx68k_bmux_1882 \mux_regs68L[7]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_2132, n_2131, n_2130, n_2129, n_2128, n_2127, n_2126,
       n_2125, n_2124, n_2123, n_2122, n_2121, n_2120, n_2119, n_2118,
       n_2117}), .z ({n_2150, n_2149, n_2148, n_2147, n_2146, n_2145,
       n_2144, n_2143, n_2142, n_2141, n_2140, n_2139, n_2138, n_2137,
       n_2136, n_2135}));
  fx68k_mux_1995 \mux_regs68L[7]_1511_27 (.ctl ({n_827, n_828}), .in_0
       (Dbd), .in_1 ({n_2150, n_2149, n_2148, n_2147, n_2146, n_2145,
       n_2144, n_2143, n_2142, n_2141, n_2140, n_2139, n_2138, n_2137,
       n_2136, n_2135}), .z ({n_2209, n_2207, n_2205, n_2203, n_2201,
       n_2199, n_2197, n_2195, n_2193, n_2191, n_2189, n_2187, n_2185,
       n_2183, n_2181, n_2179}));
  fx68k_mux_2428 \mux_regs68L[7]_1512_28 (.ctl ({n_827, n_828}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_2142, n_2141, n_2140,
       n_2139, n_2138, n_2137, n_2136, n_2135}), .z ({n_2169, n_2167,
       n_2165, n_2163, n_2161, n_2159, n_2157, n_2155}));
  fx68k_mux_1995 \mux_regs68L[7]_1513_16 (.ctl ({n_827, n_828}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_2150, n_2149, n_2148,
       n_2147, n_2146, n_2145, n_2144, n_2143, n_2142, n_2141, n_2140,
       n_2139, n_2138, n_2137, n_2136, n_2135}), .z ({n_2178, n_2177,
       n_2176, n_2175, n_2174, n_2173, n_2172, n_2171, n_2170, n_2168,
       n_2166, n_2164, n_2162, n_2160, n_2158, n_2156}));
  fx68k_bmux_1882 \mux_regs68L[7]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_2178, n_2177, n_2176, n_2175, n_2174, n_2173, n_2172,
       n_2171, n_2170, n_2168, n_2166, n_2164, n_2162, n_2160, n_2158,
       n_2156}), .in_1 ({n_2150, n_2149, n_2148, n_2147, n_2146,
       n_2145, n_2144, n_2143, n_2169, n_2167, n_2165, n_2163, n_2161,
       n_2159, n_2157, n_2155}), .z ({n_2210, n_2208, n_2206, n_2204,
       n_2202, n_2200, n_2198, n_2196, n_2194, n_2192, n_2190, n_2188,
       n_2186, n_2184, n_2182, n_2180}));
  fx68k_bmux_1882 \mux_regs68L[7]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_2210, n_2208, n_2206, n_2204, n_2202, n_2200, n_2198,
       n_2196, n_2194, n_2192, n_2190, n_2188, n_2186, n_2184, n_2182,
       n_2180}), .in_1 ({n_2209, n_2207, n_2205, n_2203, n_2201,
       n_2199, n_2197, n_2195, n_2193, n_2191, n_2189, n_2187, n_2185,
       n_2183, n_2181, n_2179}), .z ({n_2243, n_2241, n_2239, n_2237,
       n_2235, n_2233, n_2231, n_2229, n_2227, n_2225, n_2223, n_2221,
       n_2219, n_2217, n_2215, n_2213}));
  fx68k_mux_1995 \mux_regs68L[7]_1516_6 (.ctl ({n_827, n_828}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_2150, n_2149, n_2148, n_2147, n_2146,
       n_2145, n_2144, n_2143, n_2142, n_2141, n_2140, n_2139, n_2138,
       n_2137, n_2136, n_2135}), .z ({n_2244, n_2242, n_2240, n_2238,
       n_2236, n_2234, n_2232, n_2230, n_2228, n_2226, n_2224, n_2222,
       n_2220, n_2218, n_2216, n_2214}));
  fx68k_bmux_1882 \mux_regs68L[7]_1510_9 (.ctl (n_521), .in_0 ({n_2244,
       n_2242, n_2240, n_2238, n_2236, n_2234, n_2232, n_2230, n_2228,
       n_2226, n_2224, n_2222, n_2220, n_2218, n_2216, n_2214}), .in_1
       ({n_2243, n_2241, n_2239, n_2237, n_2235, n_2233, n_2231,
       n_2229, n_2227, n_2225, n_2223, n_2221, n_2219, n_2217, n_2215,
       n_2213}), .z ({n_2260, n_2259, n_2258, n_2257, n_2256, n_2255,
       n_2254, n_2253, n_2252, n_2251, n_2250, n_2249, n_2248, n_2247,
       n_2246, n_2245}));
  fx68k_bmux_1882 \mux_regs68L[7]_1509_22 (.ctl (n_520), .in_0
       ({n_2150, n_2149, n_2148, n_2147, n_2146, n_2145, n_2144,
       n_2143, n_2142, n_2141, n_2140, n_2139, n_2138, n_2137, n_2136,
       n_2135}), .in_1 ({n_2260, n_2259, n_2258, n_2257, n_2256,
       n_2255, n_2254, n_2253, n_2252, n_2251, n_2250, n_2249, n_2248,
       n_2247, n_2246, n_2245}), .z ({n_5189, n_5188, n_5187, n_5186,
       n_5185, n_5184, n_5183, n_5181, n_5180, n_5179, n_5178, n_5177,
       n_5176, n_5175, n_5174, n_5172}));
  fx68k_bmux_1882 \mux_regs68L[8]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_2276,
       n_2275, n_2274, n_2273, n_2272, n_2271, n_2270, n_2269, n_2268,
       n_2267, n_2266, n_2265, n_2264, n_2263, n_2262, n_2261}));
  fx68k_bmux_1882 \mux_regs68L[8]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_2276, n_2275, n_2274, n_2273, n_2272, n_2271, n_2270,
       n_2269, n_2268, n_2267, n_2266, n_2265, n_2264, n_2263, n_2262,
       n_2261}), .z ({n_2294, n_2293, n_2292, n_2291, n_2290, n_2289,
       n_2288, n_2287, n_2286, n_2285, n_2284, n_2283, n_2282, n_2281,
       n_2280, n_2279}));
  fx68k_mux_1995 \mux_regs68L[8]_1511_27 (.ctl ({n_845, n_846}), .in_0
       (Dbd), .in_1 ({n_2294, n_2293, n_2292, n_2291, n_2290, n_2289,
       n_2288, n_2287, n_2286, n_2285, n_2284, n_2283, n_2282, n_2281,
       n_2280, n_2279}), .z ({n_2353, n_2351, n_2349, n_2347, n_2345,
       n_2343, n_2341, n_2339, n_2337, n_2335, n_2333, n_2331, n_2329,
       n_2327, n_2325, n_2323}));
  fx68k_mux_2428 \mux_regs68L[8]_1512_28 (.ctl ({n_845, n_846}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_2286, n_2285, n_2284,
       n_2283, n_2282, n_2281, n_2280, n_2279}), .z ({n_2313, n_2311,
       n_2309, n_2307, n_2305, n_2303, n_2301, n_2299}));
  fx68k_mux_1995 \mux_regs68L[8]_1513_16 (.ctl ({n_845, n_846}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_2294, n_2293, n_2292,
       n_2291, n_2290, n_2289, n_2288, n_2287, n_2286, n_2285, n_2284,
       n_2283, n_2282, n_2281, n_2280, n_2279}), .z ({n_2322, n_2321,
       n_2320, n_2319, n_2318, n_2317, n_2316, n_2315, n_2314, n_2312,
       n_2310, n_2308, n_2306, n_2304, n_2302, n_2300}));
  fx68k_bmux_1882 \mux_regs68L[8]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_2322, n_2321, n_2320, n_2319, n_2318, n_2317, n_2316,
       n_2315, n_2314, n_2312, n_2310, n_2308, n_2306, n_2304, n_2302,
       n_2300}), .in_1 ({n_2294, n_2293, n_2292, n_2291, n_2290,
       n_2289, n_2288, n_2287, n_2313, n_2311, n_2309, n_2307, n_2305,
       n_2303, n_2301, n_2299}), .z ({n_2354, n_2352, n_2350, n_2348,
       n_2346, n_2344, n_2342, n_2340, n_2338, n_2336, n_2334, n_2332,
       n_2330, n_2328, n_2326, n_2324}));
  fx68k_bmux_1882 \mux_regs68L[8]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_2354, n_2352, n_2350, n_2348, n_2346, n_2344, n_2342,
       n_2340, n_2338, n_2336, n_2334, n_2332, n_2330, n_2328, n_2326,
       n_2324}), .in_1 ({n_2353, n_2351, n_2349, n_2347, n_2345,
       n_2343, n_2341, n_2339, n_2337, n_2335, n_2333, n_2331, n_2329,
       n_2327, n_2325, n_2323}), .z ({n_2387, n_2385, n_2383, n_2381,
       n_2379, n_2377, n_2375, n_2373, n_2371, n_2369, n_2367, n_2365,
       n_2363, n_2361, n_2359, n_2357}));
  fx68k_mux_1995 \mux_regs68L[8]_1516_6 (.ctl ({n_845, n_846}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_2294, n_2293, n_2292, n_2291, n_2290,
       n_2289, n_2288, n_2287, n_2286, n_2285, n_2284, n_2283, n_2282,
       n_2281, n_2280, n_2279}), .z ({n_2388, n_2386, n_2384, n_2382,
       n_2380, n_2378, n_2376, n_2374, n_2372, n_2370, n_2368, n_2366,
       n_2364, n_2362, n_2360, n_2358}));
  fx68k_bmux_1882 \mux_regs68L[8]_1510_9 (.ctl (n_521), .in_0 ({n_2388,
       n_2386, n_2384, n_2382, n_2380, n_2378, n_2376, n_2374, n_2372,
       n_2370, n_2368, n_2366, n_2364, n_2362, n_2360, n_2358}), .in_1
       ({n_2387, n_2385, n_2383, n_2381, n_2379, n_2377, n_2375,
       n_2373, n_2371, n_2369, n_2367, n_2365, n_2363, n_2361, n_2359,
       n_2357}), .z ({n_2404, n_2403, n_2402, n_2401, n_2400, n_2399,
       n_2398, n_2397, n_2396, n_2395, n_2394, n_2393, n_2392, n_2391,
       n_2390, n_2389}));
  fx68k_bmux_1882 \mux_regs68L[8]_1509_22 (.ctl (n_520), .in_0
       ({n_2294, n_2293, n_2292, n_2291, n_2290, n_2289, n_2288,
       n_2287, n_2286, n_2285, n_2284, n_2283, n_2282, n_2281, n_2280,
       n_2279}), .in_1 ({n_2404, n_2403, n_2402, n_2401, n_2400,
       n_2399, n_2398, n_2397, n_2396, n_2395, n_2394, n_2393, n_2392,
       n_2391, n_2390, n_2389}), .z ({n_5110, n_5109, n_5108, n_5107,
       n_5106, n_5105, n_5104, n_5102, n_5101, n_5100, n_5099, n_5098,
       n_5097, n_5096, n_5095, n_5093}));
  fx68k_bmux_1882 \mux_regs68L[9]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_2420,
       n_2419, n_2418, n_2417, n_2416, n_2415, n_2414, n_2413, n_2412,
       n_2411, n_2410, n_2409, n_2408, n_2407, n_2406, n_2405}));
  fx68k_bmux_1882 \mux_regs68L[9]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_2420, n_2419, n_2418, n_2417, n_2416, n_2415, n_2414,
       n_2413, n_2412, n_2411, n_2410, n_2409, n_2408, n_2407, n_2406,
       n_2405}), .z ({n_2438, n_2437, n_2436, n_2435, n_2434, n_2433,
       n_2432, n_2431, n_2430, n_2429, n_2428, n_2427, n_2426, n_2425,
       n_2424, n_2423}));
  fx68k_mux_1995 \mux_regs68L[9]_1511_27 (.ctl ({n_863, n_864}), .in_0
       (Dbd), .in_1 ({n_2438, n_2437, n_2436, n_2435, n_2434, n_2433,
       n_2432, n_2431, n_2430, n_2429, n_2428, n_2427, n_2426, n_2425,
       n_2424, n_2423}), .z ({n_2497, n_2495, n_2493, n_2491, n_2489,
       n_2487, n_2485, n_2483, n_2481, n_2479, n_2477, n_2475, n_2473,
       n_2471, n_2469, n_2467}));
  fx68k_mux_2428 \mux_regs68L[9]_1512_28 (.ctl ({n_863, n_864}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_2430, n_2429, n_2428,
       n_2427, n_2426, n_2425, n_2424, n_2423}), .z ({n_2457, n_2455,
       n_2453, n_2451, n_2449, n_2447, n_2445, n_2443}));
  fx68k_mux_1995 \mux_regs68L[9]_1513_16 (.ctl ({n_863, n_864}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_2438, n_2437, n_2436,
       n_2435, n_2434, n_2433, n_2432, n_2431, n_2430, n_2429, n_2428,
       n_2427, n_2426, n_2425, n_2424, n_2423}), .z ({n_2466, n_2465,
       n_2464, n_2463, n_2462, n_2461, n_2460, n_2459, n_2458, n_2456,
       n_2454, n_2452, n_2450, n_2448, n_2446, n_2444}));
  fx68k_bmux_1882 \mux_regs68L[9]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_2466, n_2465, n_2464, n_2463, n_2462, n_2461, n_2460,
       n_2459, n_2458, n_2456, n_2454, n_2452, n_2450, n_2448, n_2446,
       n_2444}), .in_1 ({n_2438, n_2437, n_2436, n_2435, n_2434,
       n_2433, n_2432, n_2431, n_2457, n_2455, n_2453, n_2451, n_2449,
       n_2447, n_2445, n_2443}), .z ({n_2498, n_2496, n_2494, n_2492,
       n_2490, n_2488, n_2486, n_2484, n_2482, n_2480, n_2478, n_2476,
       n_2474, n_2472, n_2470, n_2468}));
  fx68k_bmux_1882 \mux_regs68L[9]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_2498, n_2496, n_2494, n_2492, n_2490, n_2488, n_2486,
       n_2484, n_2482, n_2480, n_2478, n_2476, n_2474, n_2472, n_2470,
       n_2468}), .in_1 ({n_2497, n_2495, n_2493, n_2491, n_2489,
       n_2487, n_2485, n_2483, n_2481, n_2479, n_2477, n_2475, n_2473,
       n_2471, n_2469, n_2467}), .z ({n_2531, n_2529, n_2527, n_2525,
       n_2523, n_2521, n_2519, n_2517, n_2515, n_2513, n_2511, n_2509,
       n_2507, n_2505, n_2503, n_2501}));
  fx68k_mux_1995 \mux_regs68L[9]_1516_6 (.ctl ({n_863, n_864}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_2438, n_2437, n_2436, n_2435, n_2434,
       n_2433, n_2432, n_2431, n_2430, n_2429, n_2428, n_2427, n_2426,
       n_2425, n_2424, n_2423}), .z ({n_2532, n_2530, n_2528, n_2526,
       n_2524, n_2522, n_2520, n_2518, n_2516, n_2514, n_2512, n_2510,
       n_2508, n_2506, n_2504, n_2502}));
  fx68k_bmux_1882 \mux_regs68L[9]_1510_9 (.ctl (n_521), .in_0 ({n_2532,
       n_2530, n_2528, n_2526, n_2524, n_2522, n_2520, n_2518, n_2516,
       n_2514, n_2512, n_2510, n_2508, n_2506, n_2504, n_2502}), .in_1
       ({n_2531, n_2529, n_2527, n_2525, n_2523, n_2521, n_2519,
       n_2517, n_2515, n_2513, n_2511, n_2509, n_2507, n_2505, n_2503,
       n_2501}), .z ({n_2548, n_2547, n_2546, n_2545, n_2544, n_2543,
       n_2542, n_2541, n_2540, n_2539, n_2538, n_2537, n_2536, n_2535,
       n_2534, n_2533}));
  fx68k_bmux_1882 \mux_regs68L[9]_1509_22 (.ctl (n_520), .in_0
       ({n_2438, n_2437, n_2436, n_2435, n_2434, n_2433, n_2432,
       n_2431, n_2430, n_2429, n_2428, n_2427, n_2426, n_2425, n_2424,
       n_2423}), .in_1 ({n_2548, n_2547, n_2546, n_2545, n_2544,
       n_2543, n_2542, n_2541, n_2540, n_2539, n_2538, n_2537, n_2536,
       n_2535, n_2534, n_2533}), .z ({n_5031, n_5030, n_5029, n_5028,
       n_5027, n_5026, n_5025, n_5023, n_5022, n_5021, n_5020, n_5019,
       n_5018, n_5017, n_5016, n_5014}));
  fx68k_bmux_1882 \mux_regs68L[10]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_2564,
       n_2563, n_2562, n_2561, n_2560, n_2559, n_2558, n_2557, n_2556,
       n_2555, n_2554, n_2553, n_2552, n_2551, n_2550, n_2549}));
  fx68k_bmux_1882 \mux_regs68L[10]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_2564, n_2563, n_2562, n_2561, n_2560,
       n_2559, n_2558, n_2557, n_2556, n_2555, n_2554, n_2553, n_2552,
       n_2551, n_2550, n_2549}), .z ({n_2582, n_2581, n_2580, n_2579,
       n_2578, n_2577, n_2576, n_2575, n_2574, n_2573, n_2572, n_2571,
       n_2570, n_2569, n_2568, n_2567}));
  fx68k_mux_1995 \mux_regs68L[10]_1511_27 (.ctl ({n_881, n_882}), .in_0
       (Dbd), .in_1 ({n_2582, n_2581, n_2580, n_2579, n_2578, n_2577,
       n_2576, n_2575, n_2574, n_2573, n_2572, n_2571, n_2570, n_2569,
       n_2568, n_2567}), .z ({n_2641, n_2639, n_2637, n_2635, n_2633,
       n_2631, n_2629, n_2627, n_2625, n_2623, n_2621, n_2619, n_2617,
       n_2615, n_2613, n_2611}));
  fx68k_mux_2428 \mux_regs68L[10]_1512_28 (.ctl ({n_881, n_882}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_2574, n_2573, n_2572,
       n_2571, n_2570, n_2569, n_2568, n_2567}), .z ({n_2601, n_2599,
       n_2597, n_2595, n_2593, n_2591, n_2589, n_2587}));
  fx68k_mux_1995 \mux_regs68L[10]_1513_16 (.ctl ({n_881, n_882}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_2582, n_2581, n_2580,
       n_2579, n_2578, n_2577, n_2576, n_2575, n_2574, n_2573, n_2572,
       n_2571, n_2570, n_2569, n_2568, n_2567}), .z ({n_2610, n_2609,
       n_2608, n_2607, n_2606, n_2605, n_2604, n_2603, n_2602, n_2600,
       n_2598, n_2596, n_2594, n_2592, n_2590, n_2588}));
  fx68k_bmux_1882 \mux_regs68L[10]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_2610, n_2609, n_2608, n_2607, n_2606, n_2605, n_2604,
       n_2603, n_2602, n_2600, n_2598, n_2596, n_2594, n_2592, n_2590,
       n_2588}), .in_1 ({n_2582, n_2581, n_2580, n_2579, n_2578,
       n_2577, n_2576, n_2575, n_2601, n_2599, n_2597, n_2595, n_2593,
       n_2591, n_2589, n_2587}), .z ({n_2642, n_2640, n_2638, n_2636,
       n_2634, n_2632, n_2630, n_2628, n_2626, n_2624, n_2622, n_2620,
       n_2618, n_2616, n_2614, n_2612}));
  fx68k_bmux_1882 \mux_regs68L[10]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_2642, n_2640, n_2638, n_2636, n_2634, n_2632, n_2630,
       n_2628, n_2626, n_2624, n_2622, n_2620, n_2618, n_2616, n_2614,
       n_2612}), .in_1 ({n_2641, n_2639, n_2637, n_2635, n_2633,
       n_2631, n_2629, n_2627, n_2625, n_2623, n_2621, n_2619, n_2617,
       n_2615, n_2613, n_2611}), .z ({n_2675, n_2673, n_2671, n_2669,
       n_2667, n_2665, n_2663, n_2661, n_2659, n_2657, n_2655, n_2653,
       n_2651, n_2649, n_2647, n_2645}));
  fx68k_mux_1995 \mux_regs68L[10]_1516_6 (.ctl ({n_881, n_882}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_2582, n_2581, n_2580, n_2579, n_2578,
       n_2577, n_2576, n_2575, n_2574, n_2573, n_2572, n_2571, n_2570,
       n_2569, n_2568, n_2567}), .z ({n_2676, n_2674, n_2672, n_2670,
       n_2668, n_2666, n_2664, n_2662, n_2660, n_2658, n_2656, n_2654,
       n_2652, n_2650, n_2648, n_2646}));
  fx68k_bmux_1882 \mux_regs68L[10]_1510_9 (.ctl (n_521), .in_0
       ({n_2676, n_2674, n_2672, n_2670, n_2668, n_2666, n_2664,
       n_2662, n_2660, n_2658, n_2656, n_2654, n_2652, n_2650, n_2648,
       n_2646}), .in_1 ({n_2675, n_2673, n_2671, n_2669, n_2667,
       n_2665, n_2663, n_2661, n_2659, n_2657, n_2655, n_2653, n_2651,
       n_2649, n_2647, n_2645}), .z ({n_2692, n_2691, n_2690, n_2689,
       n_2688, n_2687, n_2686, n_2685, n_2684, n_2683, n_2682, n_2681,
       n_2680, n_2679, n_2678, n_2677}));
  fx68k_bmux_1882 \mux_regs68L[10]_1509_22 (.ctl (n_520), .in_0
       ({n_2582, n_2581, n_2580, n_2579, n_2578, n_2577, n_2576,
       n_2575, n_2574, n_2573, n_2572, n_2571, n_2570, n_2569, n_2568,
       n_2567}), .in_1 ({n_2692, n_2691, n_2690, n_2689, n_2688,
       n_2687, n_2686, n_2685, n_2684, n_2683, n_2682, n_2681, n_2680,
       n_2679, n_2678, n_2677}), .z ({n_4952, n_4951, n_4950, n_4949,
       n_4948, n_4947, n_4946, n_4944, n_4943, n_4942, n_4941, n_4940,
       n_4939, n_4938, n_4937, n_4935}));
  fx68k_bmux_1882 \mux_regs68L[11]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_2708,
       n_2707, n_2706, n_2705, n_2704, n_2703, n_2702, n_2701, n_2700,
       n_2699, n_2698, n_2697, n_2696, n_2695, n_2694, n_2693}));
  fx68k_bmux_1882 \mux_regs68L[11]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_2708, n_2707, n_2706, n_2705, n_2704,
       n_2703, n_2702, n_2701, n_2700, n_2699, n_2698, n_2697, n_2696,
       n_2695, n_2694, n_2693}), .z ({n_2726, n_2725, n_2724, n_2723,
       n_2722, n_2721, n_2720, n_2719, n_2718, n_2717, n_2716, n_2715,
       n_2714, n_2713, n_2712, n_2711}));
  fx68k_mux_1995 \mux_regs68L[11]_1511_27 (.ctl ({n_899, n_900}), .in_0
       (Dbd), .in_1 ({n_2726, n_2725, n_2724, n_2723, n_2722, n_2721,
       n_2720, n_2719, n_2718, n_2717, n_2716, n_2715, n_2714, n_2713,
       n_2712, n_2711}), .z ({n_2785, n_2783, n_2781, n_2779, n_2777,
       n_2775, n_2773, n_2771, n_2769, n_2767, n_2765, n_2763, n_2761,
       n_2759, n_2757, n_2755}));
  fx68k_mux_2428 \mux_regs68L[11]_1512_28 (.ctl ({n_899, n_900}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_2718, n_2717, n_2716,
       n_2715, n_2714, n_2713, n_2712, n_2711}), .z ({n_2745, n_2743,
       n_2741, n_2739, n_2737, n_2735, n_2733, n_2731}));
  fx68k_mux_1995 \mux_regs68L[11]_1513_16 (.ctl ({n_899, n_900}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_2726, n_2725, n_2724,
       n_2723, n_2722, n_2721, n_2720, n_2719, n_2718, n_2717, n_2716,
       n_2715, n_2714, n_2713, n_2712, n_2711}), .z ({n_2754, n_2753,
       n_2752, n_2751, n_2750, n_2749, n_2748, n_2747, n_2746, n_2744,
       n_2742, n_2740, n_2738, n_2736, n_2734, n_2732}));
  fx68k_bmux_1882 \mux_regs68L[11]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_2754, n_2753, n_2752, n_2751, n_2750, n_2749, n_2748,
       n_2747, n_2746, n_2744, n_2742, n_2740, n_2738, n_2736, n_2734,
       n_2732}), .in_1 ({n_2726, n_2725, n_2724, n_2723, n_2722,
       n_2721, n_2720, n_2719, n_2745, n_2743, n_2741, n_2739, n_2737,
       n_2735, n_2733, n_2731}), .z ({n_2786, n_2784, n_2782, n_2780,
       n_2778, n_2776, n_2774, n_2772, n_2770, n_2768, n_2766, n_2764,
       n_2762, n_2760, n_2758, n_2756}));
  fx68k_bmux_1882 \mux_regs68L[11]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_2786, n_2784, n_2782, n_2780, n_2778, n_2776, n_2774,
       n_2772, n_2770, n_2768, n_2766, n_2764, n_2762, n_2760, n_2758,
       n_2756}), .in_1 ({n_2785, n_2783, n_2781, n_2779, n_2777,
       n_2775, n_2773, n_2771, n_2769, n_2767, n_2765, n_2763, n_2761,
       n_2759, n_2757, n_2755}), .z ({n_2819, n_2817, n_2815, n_2813,
       n_2811, n_2809, n_2807, n_2805, n_2803, n_2801, n_2799, n_2797,
       n_2795, n_2793, n_2791, n_2789}));
  fx68k_mux_1995 \mux_regs68L[11]_1516_6 (.ctl ({n_899, n_900}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_2726, n_2725, n_2724, n_2723, n_2722,
       n_2721, n_2720, n_2719, n_2718, n_2717, n_2716, n_2715, n_2714,
       n_2713, n_2712, n_2711}), .z ({n_2820, n_2818, n_2816, n_2814,
       n_2812, n_2810, n_2808, n_2806, n_2804, n_2802, n_2800, n_2798,
       n_2796, n_2794, n_2792, n_2790}));
  fx68k_bmux_1882 \mux_regs68L[11]_1510_9 (.ctl (n_521), .in_0
       ({n_2820, n_2818, n_2816, n_2814, n_2812, n_2810, n_2808,
       n_2806, n_2804, n_2802, n_2800, n_2798, n_2796, n_2794, n_2792,
       n_2790}), .in_1 ({n_2819, n_2817, n_2815, n_2813, n_2811,
       n_2809, n_2807, n_2805, n_2803, n_2801, n_2799, n_2797, n_2795,
       n_2793, n_2791, n_2789}), .z ({n_2836, n_2835, n_2834, n_2833,
       n_2832, n_2831, n_2830, n_2829, n_2828, n_2827, n_2826, n_2825,
       n_2824, n_2823, n_2822, n_2821}));
  fx68k_bmux_1882 \mux_regs68L[11]_1509_22 (.ctl (n_520), .in_0
       ({n_2726, n_2725, n_2724, n_2723, n_2722, n_2721, n_2720,
       n_2719, n_2718, n_2717, n_2716, n_2715, n_2714, n_2713, n_2712,
       n_2711}), .in_1 ({n_2836, n_2835, n_2834, n_2833, n_2832,
       n_2831, n_2830, n_2829, n_2828, n_2827, n_2826, n_2825, n_2824,
       n_2823, n_2822, n_2821}), .z ({n_4873, n_4872, n_4871, n_4870,
       n_4869, n_4868, n_4867, n_4865, n_4864, n_4863, n_4862, n_4861,
       n_4860, n_4859, n_4858, n_4856}));
  fx68k_bmux_1882 \mux_regs68L[12]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_2852,
       n_2851, n_2850, n_2849, n_2848, n_2847, n_2846, n_2845, n_2844,
       n_2843, n_2842, n_2841, n_2840, n_2839, n_2838, n_2837}));
  fx68k_bmux_1882 \mux_regs68L[12]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_2852, n_2851, n_2850, n_2849, n_2848,
       n_2847, n_2846, n_2845, n_2844, n_2843, n_2842, n_2841, n_2840,
       n_2839, n_2838, n_2837}), .z ({n_2870, n_2869, n_2868, n_2867,
       n_2866, n_2865, n_2864, n_2863, n_2862, n_2861, n_2860, n_2859,
       n_2858, n_2857, n_2856, n_2855}));
  fx68k_mux_1995 \mux_regs68L[12]_1511_27 (.ctl ({n_917, n_918}), .in_0
       (Dbd), .in_1 ({n_2870, n_2869, n_2868, n_2867, n_2866, n_2865,
       n_2864, n_2863, n_2862, n_2861, n_2860, n_2859, n_2858, n_2857,
       n_2856, n_2855}), .z ({n_2929, n_2927, n_2925, n_2923, n_2921,
       n_2919, n_2917, n_2915, n_2913, n_2911, n_2909, n_2907, n_2905,
       n_2903, n_2901, n_2899}));
  fx68k_mux_2428 \mux_regs68L[12]_1512_28 (.ctl ({n_917, n_918}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_2862, n_2861, n_2860,
       n_2859, n_2858, n_2857, n_2856, n_2855}), .z ({n_2889, n_2887,
       n_2885, n_2883, n_2881, n_2879, n_2877, n_2875}));
  fx68k_mux_1995 \mux_regs68L[12]_1513_16 (.ctl ({n_917, n_918}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_2870, n_2869, n_2868,
       n_2867, n_2866, n_2865, n_2864, n_2863, n_2862, n_2861, n_2860,
       n_2859, n_2858, n_2857, n_2856, n_2855}), .z ({n_2898, n_2897,
       n_2896, n_2895, n_2894, n_2893, n_2892, n_2891, n_2890, n_2888,
       n_2886, n_2884, n_2882, n_2880, n_2878, n_2876}));
  fx68k_bmux_1882 \mux_regs68L[12]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_2898, n_2897, n_2896, n_2895, n_2894, n_2893, n_2892,
       n_2891, n_2890, n_2888, n_2886, n_2884, n_2882, n_2880, n_2878,
       n_2876}), .in_1 ({n_2870, n_2869, n_2868, n_2867, n_2866,
       n_2865, n_2864, n_2863, n_2889, n_2887, n_2885, n_2883, n_2881,
       n_2879, n_2877, n_2875}), .z ({n_2930, n_2928, n_2926, n_2924,
       n_2922, n_2920, n_2918, n_2916, n_2914, n_2912, n_2910, n_2908,
       n_2906, n_2904, n_2902, n_2900}));
  fx68k_bmux_1882 \mux_regs68L[12]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_2930, n_2928, n_2926, n_2924, n_2922, n_2920, n_2918,
       n_2916, n_2914, n_2912, n_2910, n_2908, n_2906, n_2904, n_2902,
       n_2900}), .in_1 ({n_2929, n_2927, n_2925, n_2923, n_2921,
       n_2919, n_2917, n_2915, n_2913, n_2911, n_2909, n_2907, n_2905,
       n_2903, n_2901, n_2899}), .z ({n_2963, n_2961, n_2959, n_2957,
       n_2955, n_2953, n_2951, n_2949, n_2947, n_2945, n_2943, n_2941,
       n_2939, n_2937, n_2935, n_2933}));
  fx68k_mux_1995 \mux_regs68L[12]_1516_6 (.ctl ({n_917, n_918}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_2870, n_2869, n_2868, n_2867, n_2866,
       n_2865, n_2864, n_2863, n_2862, n_2861, n_2860, n_2859, n_2858,
       n_2857, n_2856, n_2855}), .z ({n_2964, n_2962, n_2960, n_2958,
       n_2956, n_2954, n_2952, n_2950, n_2948, n_2946, n_2944, n_2942,
       n_2940, n_2938, n_2936, n_2934}));
  fx68k_bmux_1882 \mux_regs68L[12]_1510_9 (.ctl (n_521), .in_0
       ({n_2964, n_2962, n_2960, n_2958, n_2956, n_2954, n_2952,
       n_2950, n_2948, n_2946, n_2944, n_2942, n_2940, n_2938, n_2936,
       n_2934}), .in_1 ({n_2963, n_2961, n_2959, n_2957, n_2955,
       n_2953, n_2951, n_2949, n_2947, n_2945, n_2943, n_2941, n_2939,
       n_2937, n_2935, n_2933}), .z ({n_2980, n_2979, n_2978, n_2977,
       n_2976, n_2975, n_2974, n_2973, n_2972, n_2971, n_2970, n_2969,
       n_2968, n_2967, n_2966, n_2965}));
  fx68k_bmux_1882 \mux_regs68L[12]_1509_22 (.ctl (n_520), .in_0
       ({n_2870, n_2869, n_2868, n_2867, n_2866, n_2865, n_2864,
       n_2863, n_2862, n_2861, n_2860, n_2859, n_2858, n_2857, n_2856,
       n_2855}), .in_1 ({n_2980, n_2979, n_2978, n_2977, n_2976,
       n_2975, n_2974, n_2973, n_2972, n_2971, n_2970, n_2969, n_2968,
       n_2967, n_2966, n_2965}), .z ({n_4794, n_4793, n_4792, n_4791,
       n_4790, n_4789, n_4788, n_4786, n_4785, n_4784, n_4783, n_4782,
       n_4781, n_4780, n_4779, n_4777}));
  fx68k_bmux_1882 \mux_regs68L[13]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_2996,
       n_2995, n_2994, n_2993, n_2992, n_2991, n_2990, n_2989, n_2988,
       n_2987, n_2986, n_2985, n_2984, n_2983, n_2982, n_2981}));
  fx68k_bmux_1882 \mux_regs68L[13]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_2996, n_2995, n_2994, n_2993, n_2992,
       n_2991, n_2990, n_2989, n_2988, n_2987, n_2986, n_2985, n_2984,
       n_2983, n_2982, n_2981}), .z ({n_3014, n_3013, n_3012, n_3011,
       n_3010, n_3009, n_3008, n_3007, n_3006, n_3005, n_3004, n_3003,
       n_3002, n_3001, n_3000, n_2999}));
  fx68k_mux_1995 \mux_regs68L[13]_1511_27 (.ctl ({n_935, n_936}), .in_0
       (Dbd), .in_1 ({n_3014, n_3013, n_3012, n_3011, n_3010, n_3009,
       n_3008, n_3007, n_3006, n_3005, n_3004, n_3003, n_3002, n_3001,
       n_3000, n_2999}), .z ({n_3073, n_3071, n_3069, n_3067, n_3065,
       n_3063, n_3061, n_3059, n_3057, n_3055, n_3053, n_3051, n_3049,
       n_3047, n_3045, n_3043}));
  fx68k_mux_2428 \mux_regs68L[13]_1512_28 (.ctl ({n_935, n_936}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_3006, n_3005, n_3004,
       n_3003, n_3002, n_3001, n_3000, n_2999}), .z ({n_3033, n_3031,
       n_3029, n_3027, n_3025, n_3023, n_3021, n_3019}));
  fx68k_mux_1995 \mux_regs68L[13]_1513_16 (.ctl ({n_935, n_936}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_3014, n_3013, n_3012,
       n_3011, n_3010, n_3009, n_3008, n_3007, n_3006, n_3005, n_3004,
       n_3003, n_3002, n_3001, n_3000, n_2999}), .z ({n_3042, n_3041,
       n_3040, n_3039, n_3038, n_3037, n_3036, n_3035, n_3034, n_3032,
       n_3030, n_3028, n_3026, n_3024, n_3022, n_3020}));
  fx68k_bmux_1882 \mux_regs68L[13]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_3042, n_3041, n_3040, n_3039, n_3038, n_3037, n_3036,
       n_3035, n_3034, n_3032, n_3030, n_3028, n_3026, n_3024, n_3022,
       n_3020}), .in_1 ({n_3014, n_3013, n_3012, n_3011, n_3010,
       n_3009, n_3008, n_3007, n_3033, n_3031, n_3029, n_3027, n_3025,
       n_3023, n_3021, n_3019}), .z ({n_3074, n_3072, n_3070, n_3068,
       n_3066, n_3064, n_3062, n_3060, n_3058, n_3056, n_3054, n_3052,
       n_3050, n_3048, n_3046, n_3044}));
  fx68k_bmux_1882 \mux_regs68L[13]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_3074, n_3072, n_3070, n_3068, n_3066, n_3064, n_3062,
       n_3060, n_3058, n_3056, n_3054, n_3052, n_3050, n_3048, n_3046,
       n_3044}), .in_1 ({n_3073, n_3071, n_3069, n_3067, n_3065,
       n_3063, n_3061, n_3059, n_3057, n_3055, n_3053, n_3051, n_3049,
       n_3047, n_3045, n_3043}), .z ({n_3107, n_3105, n_3103, n_3101,
       n_3099, n_3097, n_3095, n_3093, n_3091, n_3089, n_3087, n_3085,
       n_3083, n_3081, n_3079, n_3077}));
  fx68k_mux_1995 \mux_regs68L[13]_1516_6 (.ctl ({n_935, n_936}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_3014, n_3013, n_3012, n_3011, n_3010,
       n_3009, n_3008, n_3007, n_3006, n_3005, n_3004, n_3003, n_3002,
       n_3001, n_3000, n_2999}), .z ({n_3108, n_3106, n_3104, n_3102,
       n_3100, n_3098, n_3096, n_3094, n_3092, n_3090, n_3088, n_3086,
       n_3084, n_3082, n_3080, n_3078}));
  fx68k_bmux_1882 \mux_regs68L[13]_1510_9 (.ctl (n_521), .in_0
       ({n_3108, n_3106, n_3104, n_3102, n_3100, n_3098, n_3096,
       n_3094, n_3092, n_3090, n_3088, n_3086, n_3084, n_3082, n_3080,
       n_3078}), .in_1 ({n_3107, n_3105, n_3103, n_3101, n_3099,
       n_3097, n_3095, n_3093, n_3091, n_3089, n_3087, n_3085, n_3083,
       n_3081, n_3079, n_3077}), .z ({n_3124, n_3123, n_3122, n_3121,
       n_3120, n_3119, n_3118, n_3117, n_3116, n_3115, n_3114, n_3113,
       n_3112, n_3111, n_3110, n_3109}));
  fx68k_bmux_1882 \mux_regs68L[13]_1509_22 (.ctl (n_520), .in_0
       ({n_3014, n_3013, n_3012, n_3011, n_3010, n_3009, n_3008,
       n_3007, n_3006, n_3005, n_3004, n_3003, n_3002, n_3001, n_3000,
       n_2999}), .in_1 ({n_3124, n_3123, n_3122, n_3121, n_3120,
       n_3119, n_3118, n_3117, n_3116, n_3115, n_3114, n_3113, n_3112,
       n_3111, n_3110, n_3109}), .z ({n_4715, n_4714, n_4713, n_4712,
       n_4711, n_4710, n_4709, n_4707, n_4706, n_4705, n_4704, n_4703,
       n_4702, n_4701, n_4700, n_4698}));
  fx68k_bmux_1882 \mux_regs68L[14]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_3140,
       n_3139, n_3138, n_3137, n_3136, n_3135, n_3134, n_3133, n_3132,
       n_3131, n_3130, n_3129, n_3128, n_3127, n_3126, n_3125}));
  fx68k_bmux_1882 \mux_regs68L[14]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_3140, n_3139, n_3138, n_3137, n_3136,
       n_3135, n_3134, n_3133, n_3132, n_3131, n_3130, n_3129, n_3128,
       n_3127, n_3126, n_3125}), .z ({n_3158, n_3157, n_3156, n_3155,
       n_3154, n_3153, n_3152, n_3151, n_3150, n_3149, n_3148, n_3147,
       n_3146, n_3145, n_3144, n_3143}));
  fx68k_mux_1995 \mux_regs68L[14]_1511_27 (.ctl ({n_953, n_954}), .in_0
       (Dbd), .in_1 ({n_3158, n_3157, n_3156, n_3155, n_3154, n_3153,
       n_3152, n_3151, n_3150, n_3149, n_3148, n_3147, n_3146, n_3145,
       n_3144, n_3143}), .z ({n_3217, n_3215, n_3213, n_3211, n_3209,
       n_3207, n_3205, n_3203, n_3201, n_3199, n_3197, n_3195, n_3193,
       n_3191, n_3189, n_3187}));
  fx68k_mux_2428 \mux_regs68L[14]_1512_28 (.ctl ({n_953, n_954}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_3150, n_3149, n_3148,
       n_3147, n_3146, n_3145, n_3144, n_3143}), .z ({n_3177, n_3175,
       n_3173, n_3171, n_3169, n_3167, n_3165, n_3163}));
  fx68k_mux_1995 \mux_regs68L[14]_1513_16 (.ctl ({n_953, n_954}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_3158, n_3157, n_3156,
       n_3155, n_3154, n_3153, n_3152, n_3151, n_3150, n_3149, n_3148,
       n_3147, n_3146, n_3145, n_3144, n_3143}), .z ({n_3186, n_3185,
       n_3184, n_3183, n_3182, n_3181, n_3180, n_3179, n_3178, n_3176,
       n_3174, n_3172, n_3170, n_3168, n_3166, n_3164}));
  fx68k_bmux_1882 \mux_regs68L[14]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_3186, n_3185, n_3184, n_3183, n_3182, n_3181, n_3180,
       n_3179, n_3178, n_3176, n_3174, n_3172, n_3170, n_3168, n_3166,
       n_3164}), .in_1 ({n_3158, n_3157, n_3156, n_3155, n_3154,
       n_3153, n_3152, n_3151, n_3177, n_3175, n_3173, n_3171, n_3169,
       n_3167, n_3165, n_3163}), .z ({n_3218, n_3216, n_3214, n_3212,
       n_3210, n_3208, n_3206, n_3204, n_3202, n_3200, n_3198, n_3196,
       n_3194, n_3192, n_3190, n_3188}));
  fx68k_bmux_1882 \mux_regs68L[14]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_3218, n_3216, n_3214, n_3212, n_3210, n_3208, n_3206,
       n_3204, n_3202, n_3200, n_3198, n_3196, n_3194, n_3192, n_3190,
       n_3188}), .in_1 ({n_3217, n_3215, n_3213, n_3211, n_3209,
       n_3207, n_3205, n_3203, n_3201, n_3199, n_3197, n_3195, n_3193,
       n_3191, n_3189, n_3187}), .z ({n_3251, n_3249, n_3247, n_3245,
       n_3243, n_3241, n_3239, n_3237, n_3235, n_3233, n_3231, n_3229,
       n_3227, n_3225, n_3223, n_3221}));
  fx68k_mux_1995 \mux_regs68L[14]_1516_6 (.ctl ({n_953, n_954}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_3158, n_3157, n_3156, n_3155, n_3154,
       n_3153, n_3152, n_3151, n_3150, n_3149, n_3148, n_3147, n_3146,
       n_3145, n_3144, n_3143}), .z ({n_3252, n_3250, n_3248, n_3246,
       n_3244, n_3242, n_3240, n_3238, n_3236, n_3234, n_3232, n_3230,
       n_3228, n_3226, n_3224, n_3222}));
  fx68k_bmux_1882 \mux_regs68L[14]_1510_9 (.ctl (n_521), .in_0
       ({n_3252, n_3250, n_3248, n_3246, n_3244, n_3242, n_3240,
       n_3238, n_3236, n_3234, n_3232, n_3230, n_3228, n_3226, n_3224,
       n_3222}), .in_1 ({n_3251, n_3249, n_3247, n_3245, n_3243,
       n_3241, n_3239, n_3237, n_3235, n_3233, n_3231, n_3229, n_3227,
       n_3225, n_3223, n_3221}), .z ({n_3268, n_3267, n_3266, n_3265,
       n_3264, n_3263, n_3262, n_3261, n_3260, n_3259, n_3258, n_3257,
       n_3256, n_3255, n_3254, n_3253}));
  fx68k_bmux_1882 \mux_regs68L[14]_1509_22 (.ctl (n_520), .in_0
       ({n_3158, n_3157, n_3156, n_3155, n_3154, n_3153, n_3152,
       n_3151, n_3150, n_3149, n_3148, n_3147, n_3146, n_3145, n_3144,
       n_3143}), .in_1 ({n_3268, n_3267, n_3266, n_3265, n_3264,
       n_3263, n_3262, n_3261, n_3260, n_3259, n_3258, n_3257, n_3256,
       n_3255, n_3254, n_3253}), .z ({n_4636, n_4635, n_4634, n_4633,
       n_4632, n_4631, n_4630, n_4628, n_4627, n_4626, n_4625, n_4624,
       n_4623, n_4622, n_4621, n_4619}));
  fx68k_bmux_1882 \mux_regs68L[15]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_3284,
       n_3283, n_3282, n_3281, n_3280, n_3279, n_3278, n_3277, n_3276,
       n_3275, n_3274, n_3273, n_3272, n_3271, n_3270, n_3269}));
  fx68k_bmux_1882 \mux_regs68L[15]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_3284, n_3283, n_3282, n_3281, n_3280,
       n_3279, n_3278, n_3277, n_3276, n_3275, n_3274, n_3273, n_3272,
       n_3271, n_3270, n_3269}), .z ({n_3302, n_3301, n_3300, n_3299,
       n_3298, n_3297, n_3296, n_3295, n_3294, n_3293, n_3292, n_3291,
       n_3290, n_3289, n_3288, n_3287}));
  fx68k_mux_1995 \mux_regs68L[15]_1511_27 (.ctl ({n_971, n_972}), .in_0
       (Dbd), .in_1 ({n_3302, n_3301, n_3300, n_3299, n_3298, n_3297,
       n_3296, n_3295, n_3294, n_3293, n_3292, n_3291, n_3290, n_3289,
       n_3288, n_3287}), .z ({n_3361, n_3359, n_3357, n_3355, n_3353,
       n_3351, n_3349, n_3347, n_3345, n_3343, n_3341, n_3339, n_3337,
       n_3335, n_3333, n_3331}));
  fx68k_mux_2428 \mux_regs68L[15]_1512_28 (.ctl ({n_971, n_972}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_3294, n_3293, n_3292,
       n_3291, n_3290, n_3289, n_3288, n_3287}), .z ({n_3321, n_3319,
       n_3317, n_3315, n_3313, n_3311, n_3309, n_3307}));
  fx68k_mux_1995 \mux_regs68L[15]_1513_16 (.ctl ({n_971, n_972}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_3302, n_3301, n_3300,
       n_3299, n_3298, n_3297, n_3296, n_3295, n_3294, n_3293, n_3292,
       n_3291, n_3290, n_3289, n_3288, n_3287}), .z ({n_3330, n_3329,
       n_3328, n_3327, n_3326, n_3325, n_3324, n_3323, n_3322, n_3320,
       n_3318, n_3316, n_3314, n_3312, n_3310, n_3308}));
  fx68k_bmux_1882 \mux_regs68L[15]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_3330, n_3329, n_3328, n_3327, n_3326, n_3325, n_3324,
       n_3323, n_3322, n_3320, n_3318, n_3316, n_3314, n_3312, n_3310,
       n_3308}), .in_1 ({n_3302, n_3301, n_3300, n_3299, n_3298,
       n_3297, n_3296, n_3295, n_3321, n_3319, n_3317, n_3315, n_3313,
       n_3311, n_3309, n_3307}), .z ({n_3362, n_3360, n_3358, n_3356,
       n_3354, n_3352, n_3350, n_3348, n_3346, n_3344, n_3342, n_3340,
       n_3338, n_3336, n_3334, n_3332}));
  fx68k_bmux_1882 \mux_regs68L[15]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_3362, n_3360, n_3358, n_3356, n_3354, n_3352, n_3350,
       n_3348, n_3346, n_3344, n_3342, n_3340, n_3338, n_3336, n_3334,
       n_3332}), .in_1 ({n_3361, n_3359, n_3357, n_3355, n_3353,
       n_3351, n_3349, n_3347, n_3345, n_3343, n_3341, n_3339, n_3337,
       n_3335, n_3333, n_3331}), .z ({n_3395, n_3393, n_3391, n_3389,
       n_3387, n_3385, n_3383, n_3381, n_3379, n_3377, n_3375, n_3373,
       n_3371, n_3369, n_3367, n_3365}));
  fx68k_mux_1995 \mux_regs68L[15]_1516_6 (.ctl ({n_971, n_972}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_3302, n_3301, n_3300, n_3299, n_3298,
       n_3297, n_3296, n_3295, n_3294, n_3293, n_3292, n_3291, n_3290,
       n_3289, n_3288, n_3287}), .z ({n_3396, n_3394, n_3392, n_3390,
       n_3388, n_3386, n_3384, n_3382, n_3380, n_3378, n_3376, n_3374,
       n_3372, n_3370, n_3368, n_3366}));
  fx68k_bmux_1882 \mux_regs68L[15]_1510_9 (.ctl (n_521), .in_0
       ({n_3396, n_3394, n_3392, n_3390, n_3388, n_3386, n_3384,
       n_3382, n_3380, n_3378, n_3376, n_3374, n_3372, n_3370, n_3368,
       n_3366}), .in_1 ({n_3395, n_3393, n_3391, n_3389, n_3387,
       n_3385, n_3383, n_3381, n_3379, n_3377, n_3375, n_3373, n_3371,
       n_3369, n_3367, n_3365}), .z ({n_3412, n_3411, n_3410, n_3409,
       n_3408, n_3407, n_3406, n_3405, n_3404, n_3403, n_3402, n_3401,
       n_3400, n_3399, n_3398, n_3397}));
  fx68k_bmux_1882 \mux_regs68L[15]_1509_22 (.ctl (n_520), .in_0
       ({n_3302, n_3301, n_3300, n_3299, n_3298, n_3297, n_3296,
       n_3295, n_3294, n_3293, n_3292, n_3291, n_3290, n_3289, n_3288,
       n_3287}), .in_1 ({n_3412, n_3411, n_3410, n_3409, n_3408,
       n_3407, n_3406, n_3405, n_3404, n_3403, n_3402, n_3401, n_3400,
       n_3399, n_3398, n_3397}), .z ({n_4557, n_4556, n_4555, n_4554,
       n_4553, n_4552, n_4551, n_4549, n_4548, n_4547, n_4546, n_4545,
       n_4544, n_4543, n_4542, n_4540}));
  fx68k_bmux_1882 \mux_regs68L[16]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_3428,
       n_3427, n_3426, n_3425, n_3424, n_3423, n_3422, n_3421, n_3420,
       n_3419, n_3418, n_3417, n_3416, n_3415, n_3414, n_3413}));
  fx68k_bmux_1882 \mux_regs68L[16]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_3428, n_3427, n_3426, n_3425, n_3424,
       n_3423, n_3422, n_3421, n_3420, n_3419, n_3418, n_3417, n_3416,
       n_3415, n_3414, n_3413}), .z ({n_3446, n_3445, n_3444, n_3443,
       n_3442, n_3441, n_3440, n_3439, n_3438, n_3437, n_3436, n_3435,
       n_3434, n_3433, n_3432, n_3431}));
  fx68k_mux_1995 \mux_regs68L[16]_1511_27 (.ctl ({n_989, n_990}), .in_0
       (Dbd), .in_1 ({n_3446, n_3445, n_3444, n_3443, n_3442, n_3441,
       n_3440, n_3439, n_3438, n_3437, n_3436, n_3435, n_3434, n_3433,
       n_3432, n_3431}), .z ({n_3505, n_3503, n_3501, n_3499, n_3497,
       n_3495, n_3493, n_3491, n_3489, n_3487, n_3485, n_3483, n_3481,
       n_3479, n_3477, n_3475}));
  fx68k_mux_2428 \mux_regs68L[16]_1512_28 (.ctl ({n_989, n_990}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_3438, n_3437, n_3436,
       n_3435, n_3434, n_3433, n_3432, n_3431}), .z ({n_3465, n_3463,
       n_3461, n_3459, n_3457, n_3455, n_3453, n_3451}));
  fx68k_mux_1995 \mux_regs68L[16]_1513_16 (.ctl ({n_989, n_990}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_3446, n_3445, n_3444,
       n_3443, n_3442, n_3441, n_3440, n_3439, n_3438, n_3437, n_3436,
       n_3435, n_3434, n_3433, n_3432, n_3431}), .z ({n_3474, n_3473,
       n_3472, n_3471, n_3470, n_3469, n_3468, n_3467, n_3466, n_3464,
       n_3462, n_3460, n_3458, n_3456, n_3454, n_3452}));
  fx68k_bmux_1882 \mux_regs68L[16]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_3474, n_3473, n_3472, n_3471, n_3470, n_3469, n_3468,
       n_3467, n_3466, n_3464, n_3462, n_3460, n_3458, n_3456, n_3454,
       n_3452}), .in_1 ({n_3446, n_3445, n_3444, n_3443, n_3442,
       n_3441, n_3440, n_3439, n_3465, n_3463, n_3461, n_3459, n_3457,
       n_3455, n_3453, n_3451}), .z ({n_3506, n_3504, n_3502, n_3500,
       n_3498, n_3496, n_3494, n_3492, n_3490, n_3488, n_3486, n_3484,
       n_3482, n_3480, n_3478, n_3476}));
  fx68k_bmux_1882 \mux_regs68L[16]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_3506, n_3504, n_3502, n_3500, n_3498, n_3496, n_3494,
       n_3492, n_3490, n_3488, n_3486, n_3484, n_3482, n_3480, n_3478,
       n_3476}), .in_1 ({n_3505, n_3503, n_3501, n_3499, n_3497,
       n_3495, n_3493, n_3491, n_3489, n_3487, n_3485, n_3483, n_3481,
       n_3479, n_3477, n_3475}), .z ({n_3539, n_3537, n_3535, n_3533,
       n_3531, n_3529, n_3527, n_3525, n_3523, n_3521, n_3519, n_3517,
       n_3515, n_3513, n_3511, n_3509}));
  fx68k_mux_1995 \mux_regs68L[16]_1516_6 (.ctl ({n_989, n_990}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_3446, n_3445, n_3444, n_3443, n_3442,
       n_3441, n_3440, n_3439, n_3438, n_3437, n_3436, n_3435, n_3434,
       n_3433, n_3432, n_3431}), .z ({n_3540, n_3538, n_3536, n_3534,
       n_3532, n_3530, n_3528, n_3526, n_3524, n_3522, n_3520, n_3518,
       n_3516, n_3514, n_3512, n_3510}));
  fx68k_bmux_1882 \mux_regs68L[16]_1510_9 (.ctl (n_521), .in_0
       ({n_3540, n_3538, n_3536, n_3534, n_3532, n_3530, n_3528,
       n_3526, n_3524, n_3522, n_3520, n_3518, n_3516, n_3514, n_3512,
       n_3510}), .in_1 ({n_3539, n_3537, n_3535, n_3533, n_3531,
       n_3529, n_3527, n_3525, n_3523, n_3521, n_3519, n_3517, n_3515,
       n_3513, n_3511, n_3509}), .z ({n_3556, n_3555, n_3554, n_3553,
       n_3552, n_3551, n_3550, n_3549, n_3548, n_3547, n_3546, n_3545,
       n_3544, n_3543, n_3542, n_3541}));
  fx68k_bmux_1882 \mux_regs68L[16]_1509_22 (.ctl (n_520), .in_0
       ({n_3446, n_3445, n_3444, n_3443, n_3442, n_3441, n_3440,
       n_3439, n_3438, n_3437, n_3436, n_3435, n_3434, n_3433, n_3432,
       n_3431}), .in_1 ({n_3556, n_3555, n_3554, n_3553, n_3552,
       n_3551, n_3550, n_3549, n_3548, n_3547, n_3546, n_3545, n_3544,
       n_3543, n_3542, n_3541}), .z ({n_4478, n_4477, n_4476, n_4475,
       n_4474, n_4473, n_4472, n_4470, n_4469, n_4468, n_4467, n_4466,
       n_4465, n_4464, n_4463, n_4461}));
  fx68k_bmux_1882 \mux_regs68L[17]_1501_10 (.ctl (\Nanod[dbl2rxl] ),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 (Dbd), .z ({n_3572,
       n_3571, n_3570, n_3569, n_3568, n_3567, n_3566, n_3565, n_3564,
       n_3563, n_3562, n_3561, n_3560, n_3559, n_3558, n_3557}));
  fx68k_bmux_1882 \mux_regs68L[17]_1500_9 (.ctl (n_525), .in_0
       ({n_1155, n_1153, n_1151, n_1149, n_1147, n_1145, n_1143,
       n_1141, n_1139, n_1137, n_1135, n_1133, n_1131, n_1129, n_1127,
       n_1125}), .in_1 ({n_3572, n_3571, n_3570, n_3569, n_3568,
       n_3567, n_3566, n_3565, n_3564, n_3563, n_3562, n_3561, n_3560,
       n_3559, n_3558, n_3557}), .z ({n_3590, n_3589, n_3588, n_3587,
       n_3586, n_3585, n_3584, n_3583, n_3582, n_3581, n_3580, n_3579,
       n_3578, n_3577, n_3576, n_3575}));
  fx68k_mux_1995 \mux_regs68L[17]_1511_27 (.ctl ({n_1007, n_1008}),
       .in_0 (Dbd), .in_1 ({n_3590, n_3589, n_3588, n_3587, n_3586,
       n_3585, n_3584, n_3583, n_3582, n_3581, n_3580, n_3579, n_3578,
       n_3577, n_3576, n_3575}), .z ({n_3649, n_3647, n_3645, n_3643,
       n_3641, n_3639, n_3637, n_3635, n_3633, n_3631, n_3629, n_3627,
       n_3625, n_3623, n_3621, n_3619}));
  fx68k_mux_2428 \mux_regs68L[17]_1512_28 (.ctl ({n_1007, n_1008}),
       .in_0 ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_3582, n_3581,
       n_3580, n_3579, n_3578, n_3577, n_3576, n_3575}), .z ({n_3609,
       n_3607, n_3605, n_3603, n_3601, n_3599, n_3597, n_3595}));
  fx68k_mux_1995 \mux_regs68L[17]_1513_16 (.ctl ({n_1007, n_1008}),
       .in_0 ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_3590, n_3589,
       n_3588, n_3587, n_3586, n_3585, n_3584, n_3583, n_3582, n_3581,
       n_3580, n_3579, n_3578, n_3577, n_3576, n_3575}), .z ({n_3618,
       n_3617, n_3616, n_3615, n_3614, n_3613, n_3612, n_3611, n_3610,
       n_3608, n_3606, n_3604, n_3602, n_3600, n_3598, n_3596}));
  fx68k_bmux_1882 \mux_regs68L[17]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_3618, n_3617, n_3616, n_3615, n_3614, n_3613, n_3612,
       n_3611, n_3610, n_3608, n_3606, n_3604, n_3602, n_3600, n_3598,
       n_3596}), .in_1 ({n_3590, n_3589, n_3588, n_3587, n_3586,
       n_3585, n_3584, n_3583, n_3609, n_3607, n_3605, n_3603, n_3601,
       n_3599, n_3597, n_3595}), .z ({n_3650, n_3648, n_3646, n_3644,
       n_3642, n_3640, n_3638, n_3636, n_3634, n_3632, n_3630, n_3628,
       n_3626, n_3624, n_3622, n_3620}));
  fx68k_bmux_1882 \mux_regs68L[17]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_3650, n_3648, n_3646, n_3644, n_3642, n_3640, n_3638,
       n_3636, n_3634, n_3632, n_3630, n_3628, n_3626, n_3624, n_3622,
       n_3620}), .in_1 ({n_3649, n_3647, n_3645, n_3643, n_3641,
       n_3639, n_3637, n_3635, n_3633, n_3631, n_3629, n_3627, n_3625,
       n_3623, n_3621, n_3619}), .z ({n_3683, n_3681, n_3679, n_3677,
       n_3675, n_3673, n_3671, n_3669, n_3667, n_3665, n_3663, n_3661,
       n_3659, n_3657, n_3655, n_3653}));
  fx68k_mux_1995 \mux_regs68L[17]_1516_6 (.ctl ({n_1007, n_1008}),
       .in_0 ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_3590, n_3589, n_3588, n_3587, n_3586,
       n_3585, n_3584, n_3583, n_3582, n_3581, n_3580, n_3579, n_3578,
       n_3577, n_3576, n_3575}), .z ({n_3684, n_3682, n_3680, n_3678,
       n_3676, n_3674, n_3672, n_3670, n_3668, n_3666, n_3664, n_3662,
       n_3660, n_3658, n_3656, n_3654}));
  fx68k_bmux_1882 \mux_regs68L[17]_1510_9 (.ctl (n_521), .in_0
       ({n_3684, n_3682, n_3680, n_3678, n_3676, n_3674, n_3672,
       n_3670, n_3668, n_3666, n_3664, n_3662, n_3660, n_3658, n_3656,
       n_3654}), .in_1 ({n_3683, n_3681, n_3679, n_3677, n_3675,
       n_3673, n_3671, n_3669, n_3667, n_3665, n_3663, n_3661, n_3659,
       n_3657, n_3655, n_3653}), .z ({n_3700, n_3699, n_3698, n_3697,
       n_3696, n_3695, n_3694, n_3693, n_3692, n_3691, n_3690, n_3689,
       n_3688, n_3687, n_3686, n_3685}));
  fx68k_bmux_1882 \mux_regs68L[17]_1509_22 (.ctl (n_520), .in_0
       ({n_3590, n_3589, n_3588, n_3587, n_3586, n_3585, n_3584,
       n_3583, n_3582, n_3581, n_3580, n_3579, n_3578, n_3577, n_3576,
       n_3575}), .in_1 ({n_3700, n_3699, n_3698, n_3697, n_3696,
       n_3695, n_3694, n_3693, n_3692, n_3691, n_3690, n_3689, n_3688,
       n_3687, n_3686, n_3685}), .z ({n_4399, n_4398, n_4397, n_4396,
       n_4395, n_4394, n_4393, n_4391, n_4390, n_4389, n_4388, n_4387,
       n_4386, n_4385, n_4384, n_4382}));
  fx68k_mux_2306 mux_dbdMux_1309_10(.ctl ({ryl2Dbd, rxl2Dbd,
       \Nanod[alue2Dbd] , \Nanod[dbin2Dbd] , \Nanod[alu2Dbd] ,
       \Nanod[dcr2Dbd] }), .in_0 ({\regs68L[actualRy] [15],
       \regs68L[actualRy] [14], \regs68L[actualRy] [13],
       \regs68L[actualRy] [12], \regs68L[actualRy] [11],
       \regs68L[actualRy] [10], \regs68L[actualRy] [9],
       \regs68L[actualRy] [8], \regs68L[actualRy] [7],
       \regs68L[actualRy] [6], \regs68L[actualRy] [5],
       \regs68L[actualRy] [4], \regs68L[actualRy] [3],
       \regs68L[actualRy] [2], \regs68L[actualRy] [1],
       \regs68L[actualRy] [0]}), .in_1 ({\regs68L[actualRx] [15],
       \regs68L[actualRx] [14], \regs68L[actualRx] [13],
       \regs68L[actualRx] [12], \regs68L[actualRx] [11],
       \regs68L[actualRx] [10], \regs68L[actualRx] [9],
       \regs68L[actualRx] [8], \regs68L[actualRx] [7],
       \regs68L[actualRx] [6], \regs68L[actualRx] [5],
       \regs68L[actualRx] [4], \regs68L[actualRx] [3],
       \regs68L[actualRx] [2], \regs68L[actualRx] [1],
       \regs68L[actualRx] [0]}), .in_2 (alue), .in_3 (dbin), .in_4
       (aluOut), .in_5 (dcrOutput), .z (dbdMux));
  fx68k_bmux_1503 mux_1404_18(.ctl (dblIdle), .in_0 (preDbl[15]), .in_1
       (preDbd[15]), .z (n_3766));
  fx68k_bmux_1882 mux_1406_12(.ctl (dblIdle), .in_0 (preDbl), .in_1
       (preDbd), .z ({n_3765, n_3764, n_3763, n_3762, n_3761, n_3760,
       n_3759, n_3758, n_3757, n_3756, n_3755, n_3754, n_3753, n_3752,
       n_3751, n_3750}));
  fx68k_bmux_1503 mux_1390_18(.ctl (ablIdle), .in_0 (preAbl[15]), .in_1
       (preAbd[15]), .z (n_3733));
  fx68k_bmux_1882 mux_1392_12(.ctl (ablIdle), .in_0 (preAbl), .in_1
       (preAbd), .z ({n_3732, n_3731, n_3730, n_3729, n_3728, n_3727,
       n_3726, n_3725, n_3724, n_3723, n_3722, n_3721, n_3720, n_3719,
       n_3718, n_3717}));
  fx68k_bmux_1882 mux_Abh_1391_13(.ctl (abhIdle), .in_0 (preAbh), .in_1
       ({n_3732, n_3731, n_3730, n_3729, n_3728, n_3727, n_3726,
       n_3725, n_3724, n_3723, n_3722, n_3721, n_3720, n_3719, n_3718,
       n_3717}), .z ({n_3749, n_3748, n_3747, n_3746, n_3745, n_3744,
       n_3743, n_3742, n_3741, n_3740, n_3739, n_3738, n_3737, n_3736,
       n_3735, n_3734}));
  fx68k_bmux_1882 mux_Abh_1389_8(.ctl (\Nanod[extAbh] ), .in_0
       ({n_3749, n_3748, n_3747, n_3746, n_3745, n_3744, n_3743,
       n_3742, n_3741, n_3740, n_3739, n_3738, n_3737, n_3736, n_3735,
       n_3734}), .in_1 ({n_3733, n_3733, n_3733, n_3733, n_3733,
       n_3733, n_3733, n_3733, n_3733, n_3733, n_3733, n_3733, n_3733,
       n_3733, n_3733, n_3733}), .z ({n_4242, n_4241, n_4240, n_4239,
       n_4238, n_4237, n_4236, n_4235, n_4234, n_4233, n_4232, n_4231,
       n_4230, n_4229, n_4228, n_4227}));
  fx68k_bmux_1882 mux_Dbh_1405_13(.ctl (dbhIdle), .in_0 (preDbh), .in_1
       ({n_3765, n_3764, n_3763, n_3762, n_3761, n_3760, n_3759,
       n_3758, n_3757, n_3756, n_3755, n_3754, n_3753, n_3752, n_3751,
       n_3750}), .z ({n_3782, n_3781, n_3780, n_3779, n_3778, n_3777,
       n_3776, n_3775, n_3774, n_3773, n_3772, n_3771, n_3770, n_3769,
       n_3768, n_3767}));
  fx68k_bmux_1882 mux_Dbh_1403_8(.ctl (\Nanod[extDbh] ), .in_0
       ({n_3782, n_3781, n_3780, n_3779, n_3778, n_3777, n_3776,
       n_3775, n_3774, n_3773, n_3772, n_3771, n_3770, n_3769, n_3768,
       n_3767}), .in_1 ({n_3766, n_3766, n_3766, n_3766, n_3766,
       n_3766, n_3766, n_3766, n_3766, n_3766, n_3766, n_3766, n_3766,
       n_3766, n_3766, n_3766}), .z ({n_4226, n_4225, n_4224, n_4223,
       n_4222, n_4221, n_4220, n_4219, n_4218, n_4217, n_4216, n_4215,
       n_4214, n_4213, n_4212, n_4211}));
  fx68k_bmux_1882 mux_1399_12(.ctl (\Nanod[ablAbh] ), .in_0 (preAbd),
       .in_1 (preAbh), .z ({n_3798, n_3797, n_3796, n_3795, n_3794,
       n_3793, n_3792, n_3791, n_3790, n_3789, n_3788, n_3787, n_3786,
       n_3785, n_3784, n_3783}));
  fx68k_bmux_1882 mux_Abl_1396_8(.ctl (n_552), .in_0 ({n_3798, n_3797,
       n_3796, n_3795, n_3794, n_3793, n_3792, n_3791, n_3790, n_3789,
       n_3788, n_3787, n_3786, n_3785, n_3784, n_3783}), .in_1
       (preAbl), .z (Abl));
  fx68k_bmux_1882 \mux_regs68L[1]_1500_9 (.ctl (n_525), .in_0 ({n_1155,
       n_1153, n_1151, n_1149, n_1147, n_1145, n_1143, n_1141, n_1139,
       n_1137, n_1135, n_1133, n_1131, n_1129, n_1127, n_1125}), .in_1
       ({n_3814, n_3813, n_3812, n_3811, n_3810, n_3809, n_3808,
       n_3807, n_3806, n_3805, n_3804, n_3803, n_3802, n_3801, n_3800,
       n_3799}), .z ({n_3832, n_3831, n_3830, n_3829, n_3828, n_3827,
       n_3826, n_3825, n_3824, n_3823, n_3822, n_3821, n_3820, n_3819,
       n_3818, n_3817}));
  fx68k_mux_1995 \mux_regs68L[1]_1511_27 (.ctl ({n_719, n_720}), .in_0
       (Dbd), .in_1 ({n_3832, n_3831, n_3830, n_3829, n_3828, n_3827,
       n_3826, n_3825, n_3824, n_3823, n_3822, n_3821, n_3820, n_3819,
       n_3818, n_3817}), .z ({n_3891, n_3889, n_3887, n_3885, n_3883,
       n_3881, n_3879, n_3877, n_3875, n_3873, n_3871, n_3869, n_3867,
       n_3865, n_3863, n_3861}));
  fx68k_mux_2428 \mux_regs68L[1]_1512_28 (.ctl ({n_719, n_720}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_3824, n_3823, n_3822,
       n_3821, n_3820, n_3819, n_3818, n_3817}), .z ({n_3851, n_3849,
       n_3847, n_3845, n_3843, n_3841, n_3839, n_3837}));
  fx68k_mux_1995 \mux_regs68L[1]_1513_16 (.ctl ({n_719, n_720}), .in_0
       ({Abd[15:3], dcrInput[2:0]}), .in_1 ({n_3832, n_3831, n_3830,
       n_3829, n_3828, n_3827, n_3826, n_3825, n_3824, n_3823, n_3822,
       n_3821, n_3820, n_3819, n_3818, n_3817}), .z ({n_3860, n_3859,
       n_3858, n_3857, n_3856, n_3855, n_3854, n_3853, n_3852, n_3850,
       n_3848, n_3846, n_3844, n_3842, n_3840, n_3838}));
  fx68k_bmux_1882 \mux_regs68L[1]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_3860, n_3859, n_3858, n_3857, n_3856, n_3855, n_3854,
       n_3853, n_3852, n_3850, n_3848, n_3846, n_3844, n_3842, n_3840,
       n_3838}), .in_1 ({n_3832, n_3831, n_3830, n_3829, n_3828,
       n_3827, n_3826, n_3825, n_3851, n_3849, n_3847, n_3845, n_3843,
       n_3841, n_3839, n_3837}), .z ({n_3892, n_3890, n_3888, n_3886,
       n_3884, n_3882, n_3880, n_3878, n_3876, n_3874, n_3872, n_3870,
       n_3868, n_3866, n_3864, n_3862}));
  fx68k_bmux_1882 \mux_regs68L[1]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_3892, n_3890, n_3888, n_3886, n_3884, n_3882, n_3880,
       n_3878, n_3876, n_3874, n_3872, n_3870, n_3868, n_3866, n_3864,
       n_3862}), .in_1 ({n_3891, n_3889, n_3887, n_3885, n_3883,
       n_3881, n_3879, n_3877, n_3875, n_3873, n_3871, n_3869, n_3867,
       n_3865, n_3863, n_3861}), .z ({n_3925, n_3923, n_3921, n_3919,
       n_3917, n_3915, n_3913, n_3911, n_3909, n_3907, n_3905, n_3903,
       n_3901, n_3899, n_3897, n_3895}));
  fx68k_mux_1995 \mux_regs68L[1]_1516_6 (.ctl ({n_719, n_720}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_3832, n_3831, n_3830, n_3829, n_3828,
       n_3827, n_3826, n_3825, n_3824, n_3823, n_3822, n_3821, n_3820,
       n_3819, n_3818, n_3817}), .z ({n_3926, n_3924, n_3922, n_3920,
       n_3918, n_3916, n_3914, n_3912, n_3910, n_3908, n_3906, n_3904,
       n_3902, n_3900, n_3898, n_3896}));
  fx68k_bmux_1882 \mux_regs68L[1]_1510_9 (.ctl (n_521), .in_0 ({n_3926,
       n_3924, n_3922, n_3920, n_3918, n_3916, n_3914, n_3912, n_3910,
       n_3908, n_3906, n_3904, n_3902, n_3900, n_3898, n_3896}), .in_1
       ({n_3925, n_3923, n_3921, n_3919, n_3917, n_3915, n_3913,
       n_3911, n_3909, n_3907, n_3905, n_3903, n_3901, n_3899, n_3897,
       n_3895}), .z ({n_3942, n_3941, n_3940, n_3939, n_3938, n_3937,
       n_3936, n_3935, n_3934, n_3933, n_3932, n_3931, n_3930, n_3929,
       n_3928, n_3927}));
  fx68k_bmux_1882 \mux_regs68L[1]_1509_22 (.ctl (n_520), .in_0
       ({n_3832, n_3831, n_3830, n_3829, n_3828, n_3827, n_3826,
       n_3825, n_3824, n_3823, n_3822, n_3821, n_3820, n_3819, n_3818,
       n_3817}), .in_1 ({n_3942, n_3941, n_3940, n_3939, n_3938,
       n_3937, n_3936, n_3935, n_3934, n_3933, n_3932, n_3931, n_3930,
       n_3929, n_3928, n_3927}), .z ({n_5663, n_5662, n_5661, n_5660,
       n_5659, n_5658, n_5657, n_5655, n_5654, n_5653, n_5652, n_5651,
       n_5650, n_5649, n_5648, n_5646}));
  fx68k_mux_2428 \mux_regs68L[0]_1512_28 (.ctl ({n_669, n_670}), .in_0
       ({Abd[7:3], dcrInput[2:0]}), .in_1 ({n_1165, n_1164, n_1163,
       n_1162, n_1161, n_1160, n_1159, n_1158}), .z ({n_3959, n_3957,
       n_3955, n_3953, n_3951, n_3949, n_3947, n_3945}));
  fx68k_bmux_1882 \mux_regs68L[0]_1512_15 (.ctl (abdIsByte), .in_0
       ({n_3968, n_3967, n_3966, n_3965, n_3964, n_3963, n_3962,
       n_3961, n_3960, n_3958, n_3956, n_3954, n_3952, n_3950, n_3948,
       n_3946}), .in_1 ({n_1173, n_1172, n_1171, n_1170, n_1169,
       n_1168, n_1167, n_1166, n_3959, n_3957, n_3955, n_3953, n_3951,
       n_3949, n_3947, n_3945}), .z ({n_4000, n_3998, n_3996, n_3994,
       n_3992, n_3990, n_3988, n_3986, n_3984, n_3982, n_3980, n_3978,
       n_3976, n_3974, n_3972, n_3970}));
  fx68k_bmux_1882 \mux_regs68L[0]_1511_10 (.ctl (\Nanod[dbl2ryl] ),
       .in_0 ({n_4000, n_3998, n_3996, n_3994, n_3992, n_3990, n_3988,
       n_3986, n_3984, n_3982, n_3980, n_3978, n_3976, n_3974, n_3972,
       n_3970}), .in_1 ({n_3999, n_3997, n_3995, n_3993, n_3991,
       n_3989, n_3987, n_3985, n_3983, n_3981, n_3979, n_3977, n_3975,
       n_3973, n_3971, n_3969}), .z ({n_4033, n_4031, n_4029, n_4027,
       n_4025, n_4023, n_4021, n_4019, n_4017, n_4015, n_4013, n_4011,
       n_4009, n_4007, n_4005, n_4003}));
  fx68k_mux_1995 \mux_regs68L[0]_1516_6 (.ctl ({n_669, n_670}), .in_0
       ({n_1492, n_1491, n_1490, n_1489, n_1488, n_1487, n_1486,
       n_1485, n_1484, n_1483, n_1482, n_1481, n_1480, n_1479, n_1478,
       n_1477}), .in_1 ({n_1173, n_1172, n_1171, n_1170, n_1169,
       n_1168, n_1167, n_1166, n_1165, n_1164, n_1163, n_1162, n_1161,
       n_1160, n_1159, n_1158}), .z ({n_4034, n_4032, n_4030, n_4028,
       n_4026, n_4024, n_4022, n_4020, n_4018, n_4016, n_4014, n_4012,
       n_4010, n_4008, n_4006, n_4004}));
  fx68k_bmux_1882 \mux_regs68L[0]_1510_9 (.ctl (n_521), .in_0 ({n_4034,
       n_4032, n_4030, n_4028, n_4026, n_4024, n_4022, n_4020, n_4018,
       n_4016, n_4014, n_4012, n_4010, n_4008, n_4006, n_4004}), .in_1
       ({n_4033, n_4031, n_4029, n_4027, n_4025, n_4023, n_4021,
       n_4019, n_4017, n_4015, n_4013, n_4011, n_4009, n_4007, n_4005,
       n_4003}), .z ({n_4050, n_4049, n_4048, n_4047, n_4046, n_4045,
       n_4044, n_4043, n_4042, n_4041, n_4040, n_4039, n_4038, n_4037,
       n_4036, n_4035}));
  fx68k_bmux_1882 \mux_regs68L[0]_1509_22 (.ctl (n_520), .in_0
       ({n_1173, n_1172, n_1171, n_1170, n_1169, n_1168, n_1167,
       n_1166, n_1165, n_1164, n_1163, n_1162, n_1161, n_1160, n_1159,
       n_1158}), .in_1 ({n_4050, n_4049, n_4048, n_4047, n_4046,
       n_4045, n_4044, n_4043, n_4042, n_4041, n_4040, n_4039, n_4038,
       n_4037, n_4036, n_4035}), .z ({n_5742, n_5741, n_5740, n_5739,
       n_5738, n_5737, n_5736, n_5734, n_5733, n_5732, n_5731, n_5730,
       n_5729, n_5728, n_5727, n_5725}));
  fx68k_bmux_1503 mux_1275_41(.ctl (\Nanod[rxlDbl] ), .in_0 (ryIsSp),
       .in_1 (rxIsSp), .z (n_4181));
  and g3 (n_8, \Irdecod[rxIsDt] , n_4178);
  and g6 (n_449, \Irdecod[ryIsDt] , n_4179);
  and g8 (n_523, n_1344, pswS);
  not g9 (n_4182, n_4181);
  and g10 (n_4184, \Irdecod[isByte] , n_4182);
  or g11 (n_4185, rxIsSp, rxMux[3]);
  or g12 (n_4186, ryIsSp, ryMux[3]);
  and g13 (n_4183, \Nanod[abdIsByte] , \Irdecod[isByte] );
  or g20 (n_4187, ryIsAreg, \Nanod[ablAbd] );
  and g21 (ryl2Abl, \Nanod[ryl2ab] , n_4187);
  not g22 (n_521, ryIsAreg);
  or g23 (n_4188, n_521, \Nanod[ablAbd] );
  and g24 (ryl2Abd, \Nanod[ryl2ab] , n_4188);
  or g25 (n_4189, ryIsAreg, \Nanod[dblDbd] );
  and g26 (ryl2Dbl, \Nanod[ryl2db] , n_4189);
  or g27 (n_4190, n_521, \Nanod[dblDbd] );
  and g28 (ryl2Dbd, \Nanod[ryl2db] , n_4190);
  or g29 (n_4191, rxIsAreg, \Nanod[ablAbd] );
  and g30 (rxl2Abl, \Nanod[rxl2ab] , n_4191);
  not g31 (n_525, rxIsAreg);
  or g32 (n_4192, n_525, \Nanod[ablAbd] );
  and g33 (rxl2Abd, \Nanod[rxl2ab] , n_4192);
  or g34 (n_4193, rxIsAreg, \Nanod[dblDbd] );
  and g35 (rxl2Dbl, \Nanod[rxl2db] , n_4193);
  or g36 (n_4194, n_525, \Nanod[dblDbd] );
  and g37 (rxl2Dbd, \Nanod[rxl2db] , n_4194);
  not g38 (n_552, ablIdle);
  not g39 (n_536, abdIdle);
  not g40 (n_518, dblIdle);
  not g41 (n_1358, dbdIdle);
  and g54 (n_4275, \Nanod[au2Db] , \Nanod[db2Aob] );
  or g55 (au2Aob, \Nanod[au2Aob] , n_4275);
  and g56 (n_451, enT1, au2Aob);
  or g60 (n_1226, byteNotSpAlign, \Nanod[noSpAlign] );
  and g62 (n_453, enT3, \Nanod[auClkEn] );
  or g64 (n_524, \Nanod[dbl2rxl] , \Nanod[abl2rxl] );
  or g65 (n_520, \Nanod[dbl2ryl] , \Nanod[abl2ryl] );
  or g66 (n_667, \Nanod[dbh2rxh] , \Nanod[abh2rxh] );
  or g67 (n_654, \Nanod[dbh2ryh] , \Nanod[abh2ryh] );
  and g104 (n_554, \Nanod[dbl2reg] , \Nanod[pcldbl] );
  and g105 (n_641, \Nanod[dbh2reg] , \Nanod[pchdbh] );
  and g106 (n_1027, \Nanod[abh2reg] , \Nanod[pchabh] );
  and g107 (n_555, \Nanod[abl2reg] , \Nanod[pclabl] );
  and g108 (n_505, \Nanod[reg2dbl] , \Nanod[pcldbl] );
  and g109 (n_644, \Nanod[reg2dbh] , \Nanod[pchdbh] );
  and g110 (n_537, \Nanod[reg2abl] , \Nanod[pclabl] );
  and g111 (n_639, \Nanod[reg2abh] , \Nanod[pchabh] );
  and g112 (n_553, enT1, \Nanod[au2Pc] );
  and g127 (n_456, enT1, \Nanod[abl2Pren] );
  and g128 (n_457, enT3, \Nanod[updPren] );
  and g147 (n_643, enT3, \Nanod[abd2Dcr] );
  and g151 (alueClkEn, enT3, \Nanod[dbd2Alue] );
  not g157 (n_6288, \Nanod[dbd2Alub] );
  not g162 (n_4280, n_451);
  not g163 (n_6286, \Clks[pwrUp] );
  not g167 (n_6262, n_456);
  not g174 (n_4375, n_520);
  not g176 (n_4356, \Nanod[dbl2ryl] );
  not g180 (n_4322, \Nanod[dbl2rxl] );
  not g181 (n_4318, abdIsByte);
  not g184 (n_6180, n_553);
  not g185 (n_6176, dbl2Pcl);
  not g187 (n_6242, \Nanod[dbl2Atl] );
  not g191 (n_6199, dbh2Pch);
  not g196 (n_5747, n_654);
  not g203 (n_670, n_669);
  not g204 (n_720, n_719);
  not g205 (n_738, n_737);
  not g206 (n_756, n_755);
  not g207 (n_774, n_773);
  not g208 (n_792, n_791);
  not g209 (n_810, n_809);
  not g210 (n_828, n_827);
  not g211 (n_846, n_845);
  not g212 (n_864, n_863);
  not g213 (n_882, n_881);
  not g214 (n_900, n_899);
  not g215 (n_918, n_917);
  not g216 (n_936, n_935);
  not g217 (n_954, n_953);
  not g218 (n_972, n_971);
  not g219 (n_990, n_989);
  not g220 (n_1008, n_1007);
  not g221 (n_6222, \Nanod[abh2Ath] );
  not g230 (n_4276, \Nanod[db2Aob] );
  CDN_dc logicX_inst(.cf (1'b0), .dcf (1'b1), .z (_X_));
  and g306 (n_4277, \Nanod[ab2Aob] , n_4276);
  or g307 (n_4278, n_4277, \Nanod[db2Aob] );
  and g308 (n_4279, n_4278, enT2);
  and g309 (n_4281, n_4279, n_4280);
  or g310 (n_4283, n_4281, n_451);
  and g311 (n_4324, n_4315, \Nanod[dbl2rxl] );
  and g312 (n_4320, n_4315, abdIsByte);
  and g313 (n_4319, n_4315, n_4318);
  or g314 (n_4321, n_4319, n_4320);
  and g316 (n_4323, n_4321, n_4322);
  or g317 (n_4327, n_4323, n_4324);
  and g318 (n_4326, n_4319, n_4322);
  or g319 (n_4328, n_4326, n_4324);
  and g320 (n_4332, n_4327, n_525);
  and g321 (n_4334, n_4328, n_525);
  and g322 (n_4331, n_4315, rxIsAreg);
  or g323 (n_4335, n_4331, n_4332);
  or g325 (n_4336, n_4331, n_4334);
  and g326 (n_4337, n_4335, n_524);
  and g327 (n_4339, n_4336, n_524);
  and g328 (n_4338, n_4337, n_1008);
  or g329 (n_4341, n_4338, n_1007);
  and g330 (n_4340, n_4339, n_1008);
  or g331 (n_4342, n_4340, n_1007);
  and g332 (n_4358, n_4341, \Nanod[dbl2ryl] );
  and g333 (n_4361, n_4342, \Nanod[dbl2ryl] );
  and g339 (n_4351, n_4341, abdIsByte);
  and g340 (n_4354, n_4339, abdIsByte);
  and g345 (n_4350, n_4341, n_4318);
  or g346 (n_4355, n_4350, n_4351);
  and g347 (n_4353, n_4342, n_4318);
  or g348 (n_4359, n_4353, n_4354);
  and g349 (n_4357, n_4355, n_4356);
  or g350 (n_4362, n_4357, n_4358);
  and g351 (n_4360, n_4359, n_4356);
  or g352 (n_4363, n_4360, n_4361);
  and g353 (n_4369, n_4362, n_521);
  and g354 (n_4372, n_4363, n_521);
  and g359 (n_4368, n_4341, ryIsAreg);
  or g360 (n_4373, n_4368, n_4369);
  and g361 (n_4371, n_4342, ryIsAreg);
  or g362 (n_4374, n_4371, n_4372);
  and g363 (n_4377, n_4373, n_520);
  and g364 (n_4379, n_4374, n_520);
  and g365 (n_4376, n_4337, n_4375);
  or g366 (n_4380, n_4376, n_4377);
  and g367 (n_4378, n_4339, n_4375);
  or g368 (n_4381, n_4378, n_4379);
  and g369 (n_4383, n_4380, enT3);
  and g370 (n_4392, n_4381, enT3);
  and g371 (n_4407, n_4400, \Nanod[dbl2rxl] );
  and g372 (n_4404, n_4400, abdIsByte);
  and g373 (n_4403, n_4400, n_4318);
  or g374 (n_4405, n_4403, n_4404);
  and g376 (n_4406, n_4405, n_4322);
  or g377 (n_4410, n_4406, n_4407);
  and g378 (n_4409, n_4403, n_4322);
  or g379 (n_4411, n_4409, n_4407);
  and g380 (n_4414, n_4410, n_525);
  and g381 (n_4416, n_4411, n_525);
  and g382 (n_4413, n_4400, rxIsAreg);
  or g383 (n_4417, n_4413, n_4414);
  or g385 (n_4418, n_4413, n_4416);
  and g386 (n_4419, n_4417, n_524);
  and g387 (n_4421, n_4418, n_524);
  and g388 (n_4420, n_4419, n_990);
  or g389 (n_4423, n_4420, n_989);
  and g390 (n_4422, n_4421, n_990);
  or g391 (n_4424, n_4422, n_989);
  and g392 (n_4439, n_4423, \Nanod[dbl2ryl] );
  and g393 (n_4442, n_4424, \Nanod[dbl2ryl] );
  and g399 (n_4433, n_4423, abdIsByte);
  and g400 (n_4436, n_4421, abdIsByte);
  and g405 (n_4432, n_4423, n_4318);
  or g406 (n_4437, n_4432, n_4433);
  and g407 (n_4435, n_4424, n_4318);
  or g408 (n_4440, n_4435, n_4436);
  and g409 (n_4438, n_4437, n_4356);
  or g410 (n_4443, n_4438, n_4439);
  and g411 (n_4441, n_4440, n_4356);
  or g412 (n_4444, n_4441, n_4442);
  and g413 (n_4449, n_4443, n_521);
  and g414 (n_4452, n_4444, n_521);
  and g419 (n_4448, n_4423, ryIsAreg);
  or g420 (n_4453, n_4448, n_4449);
  and g421 (n_4451, n_4424, ryIsAreg);
  or g422 (n_4454, n_4451, n_4452);
  and g423 (n_4456, n_4453, n_520);
  and g424 (n_4458, n_4454, n_520);
  and g425 (n_4455, n_4419, n_4375);
  or g426 (n_4459, n_4455, n_4456);
  and g427 (n_4457, n_4421, n_4375);
  or g428 (n_4460, n_4457, n_4458);
  and g429 (n_4462, n_4459, enT3);
  and g430 (n_4471, n_4460, enT3);
  and g431 (n_4486, n_4479, \Nanod[dbl2rxl] );
  and g432 (n_4483, n_4479, abdIsByte);
  and g433 (n_4482, n_4479, n_4318);
  or g434 (n_4484, n_4482, n_4483);
  and g436 (n_4485, n_4484, n_4322);
  or g437 (n_4489, n_4485, n_4486);
  and g438 (n_4488, n_4482, n_4322);
  or g439 (n_4490, n_4488, n_4486);
  and g440 (n_4493, n_4489, n_525);
  and g441 (n_4495, n_4490, n_525);
  and g442 (n_4492, n_4479, rxIsAreg);
  or g443 (n_4496, n_4492, n_4493);
  or g445 (n_4497, n_4492, n_4495);
  and g446 (n_4498, n_4496, n_524);
  and g447 (n_4500, n_4497, n_524);
  and g448 (n_4499, n_4498, n_972);
  or g449 (n_4502, n_4499, n_971);
  and g450 (n_4501, n_4500, n_972);
  or g451 (n_4503, n_4501, n_971);
  and g452 (n_4518, n_4502, \Nanod[dbl2ryl] );
  and g453 (n_4521, n_4503, \Nanod[dbl2ryl] );
  and g459 (n_4512, n_4502, abdIsByte);
  and g460 (n_4515, n_4500, abdIsByte);
  and g465 (n_4511, n_4502, n_4318);
  or g466 (n_4516, n_4511, n_4512);
  and g467 (n_4514, n_4503, n_4318);
  or g468 (n_4519, n_4514, n_4515);
  and g469 (n_4517, n_4516, n_4356);
  or g470 (n_4522, n_4517, n_4518);
  and g471 (n_4520, n_4519, n_4356);
  or g472 (n_4523, n_4520, n_4521);
  and g473 (n_4528, n_4522, n_521);
  and g474 (n_4531, n_4523, n_521);
  and g479 (n_4527, n_4502, ryIsAreg);
  or g480 (n_4532, n_4527, n_4528);
  and g481 (n_4530, n_4503, ryIsAreg);
  or g482 (n_4533, n_4530, n_4531);
  and g483 (n_4535, n_4532, n_520);
  and g484 (n_4537, n_4533, n_520);
  and g485 (n_4534, n_4498, n_4375);
  or g486 (n_4538, n_4534, n_4535);
  and g487 (n_4536, n_4500, n_4375);
  or g488 (n_4539, n_4536, n_4537);
  and g489 (n_4541, n_4538, enT3);
  and g490 (n_4550, n_4539, enT3);
  and g491 (n_4565, n_4558, \Nanod[dbl2rxl] );
  and g492 (n_4562, n_4558, abdIsByte);
  and g493 (n_4561, n_4558, n_4318);
  or g494 (n_4563, n_4561, n_4562);
  and g496 (n_4564, n_4563, n_4322);
  or g497 (n_4568, n_4564, n_4565);
  and g498 (n_4567, n_4561, n_4322);
  or g499 (n_4569, n_4567, n_4565);
  and g500 (n_4572, n_4568, n_525);
  and g501 (n_4574, n_4569, n_525);
  and g502 (n_4571, n_4558, rxIsAreg);
  or g503 (n_4575, n_4571, n_4572);
  or g505 (n_4576, n_4571, n_4574);
  and g506 (n_4577, n_4575, n_524);
  and g507 (n_4579, n_4576, n_524);
  and g508 (n_4578, n_4577, n_954);
  or g509 (n_4581, n_4578, n_953);
  and g510 (n_4580, n_4579, n_954);
  or g511 (n_4582, n_4580, n_953);
  and g512 (n_4597, n_4581, \Nanod[dbl2ryl] );
  and g513 (n_4600, n_4582, \Nanod[dbl2ryl] );
  and g519 (n_4591, n_4581, abdIsByte);
  and g520 (n_4594, n_4579, abdIsByte);
  and g525 (n_4590, n_4581, n_4318);
  or g526 (n_4595, n_4590, n_4591);
  and g527 (n_4593, n_4582, n_4318);
  or g528 (n_4598, n_4593, n_4594);
  and g529 (n_4596, n_4595, n_4356);
  or g530 (n_4601, n_4596, n_4597);
  and g531 (n_4599, n_4598, n_4356);
  or g532 (n_4602, n_4599, n_4600);
  and g533 (n_4607, n_4601, n_521);
  and g534 (n_4610, n_4602, n_521);
  and g539 (n_4606, n_4581, ryIsAreg);
  or g540 (n_4611, n_4606, n_4607);
  and g541 (n_4609, n_4582, ryIsAreg);
  or g542 (n_4612, n_4609, n_4610);
  and g543 (n_4614, n_4611, n_520);
  and g544 (n_4616, n_4612, n_520);
  and g545 (n_4613, n_4577, n_4375);
  or g546 (n_4617, n_4613, n_4614);
  and g547 (n_4615, n_4579, n_4375);
  or g548 (n_4618, n_4615, n_4616);
  and g549 (n_4620, n_4617, enT3);
  and g550 (n_4629, n_4618, enT3);
  and g551 (n_4644, n_4637, \Nanod[dbl2rxl] );
  and g552 (n_4641, n_4637, abdIsByte);
  and g553 (n_4640, n_4637, n_4318);
  or g554 (n_4642, n_4640, n_4641);
  and g556 (n_4643, n_4642, n_4322);
  or g557 (n_4647, n_4643, n_4644);
  and g558 (n_4646, n_4640, n_4322);
  or g559 (n_4648, n_4646, n_4644);
  and g560 (n_4651, n_4647, n_525);
  and g561 (n_4653, n_4648, n_525);
  and g562 (n_4650, n_4637, rxIsAreg);
  or g563 (n_4654, n_4650, n_4651);
  or g565 (n_4655, n_4650, n_4653);
  and g566 (n_4656, n_4654, n_524);
  and g567 (n_4658, n_4655, n_524);
  and g568 (n_4657, n_4656, n_936);
  or g569 (n_4660, n_4657, n_935);
  and g570 (n_4659, n_4658, n_936);
  or g571 (n_4661, n_4659, n_935);
  and g572 (n_4676, n_4660, \Nanod[dbl2ryl] );
  and g573 (n_4679, n_4661, \Nanod[dbl2ryl] );
  and g579 (n_4670, n_4660, abdIsByte);
  and g580 (n_4673, n_4658, abdIsByte);
  and g585 (n_4669, n_4660, n_4318);
  or g586 (n_4674, n_4669, n_4670);
  and g587 (n_4672, n_4661, n_4318);
  or g588 (n_4677, n_4672, n_4673);
  and g589 (n_4675, n_4674, n_4356);
  or g590 (n_4680, n_4675, n_4676);
  and g591 (n_4678, n_4677, n_4356);
  or g592 (n_4681, n_4678, n_4679);
  and g593 (n_4686, n_4680, n_521);
  and g594 (n_4689, n_4681, n_521);
  and g599 (n_4685, n_4660, ryIsAreg);
  or g600 (n_4690, n_4685, n_4686);
  and g601 (n_4688, n_4661, ryIsAreg);
  or g602 (n_4691, n_4688, n_4689);
  and g603 (n_4693, n_4690, n_520);
  and g604 (n_4695, n_4691, n_520);
  and g605 (n_4692, n_4656, n_4375);
  or g606 (n_4696, n_4692, n_4693);
  and g607 (n_4694, n_4658, n_4375);
  or g608 (n_4697, n_4694, n_4695);
  and g609 (n_4699, n_4696, enT3);
  and g610 (n_4708, n_4697, enT3);
  and g611 (n_4723, n_4716, \Nanod[dbl2rxl] );
  and g612 (n_4720, n_4716, abdIsByte);
  and g613 (n_4719, n_4716, n_4318);
  or g614 (n_4721, n_4719, n_4720);
  and g616 (n_4722, n_4721, n_4322);
  or g617 (n_4726, n_4722, n_4723);
  and g618 (n_4725, n_4719, n_4322);
  or g619 (n_4727, n_4725, n_4723);
  and g620 (n_4730, n_4726, n_525);
  and g621 (n_4732, n_4727, n_525);
  and g622 (n_4729, n_4716, rxIsAreg);
  or g623 (n_4733, n_4729, n_4730);
  or g625 (n_4734, n_4729, n_4732);
  and g626 (n_4735, n_4733, n_524);
  and g627 (n_4737, n_4734, n_524);
  and g628 (n_4736, n_4735, n_918);
  or g629 (n_4739, n_4736, n_917);
  and g630 (n_4738, n_4737, n_918);
  or g631 (n_4740, n_4738, n_917);
  and g632 (n_4755, n_4739, \Nanod[dbl2ryl] );
  and g633 (n_4758, n_4740, \Nanod[dbl2ryl] );
  and g639 (n_4749, n_4739, abdIsByte);
  and g640 (n_4752, n_4737, abdIsByte);
  and g645 (n_4748, n_4739, n_4318);
  or g646 (n_4753, n_4748, n_4749);
  and g647 (n_4751, n_4740, n_4318);
  or g648 (n_4756, n_4751, n_4752);
  and g649 (n_4754, n_4753, n_4356);
  or g650 (n_4759, n_4754, n_4755);
  and g651 (n_4757, n_4756, n_4356);
  or g652 (n_4760, n_4757, n_4758);
  and g653 (n_4765, n_4759, n_521);
  and g654 (n_4768, n_4760, n_521);
  and g659 (n_4764, n_4739, ryIsAreg);
  or g660 (n_4769, n_4764, n_4765);
  and g661 (n_4767, n_4740, ryIsAreg);
  or g662 (n_4770, n_4767, n_4768);
  and g663 (n_4772, n_4769, n_520);
  and g664 (n_4774, n_4770, n_520);
  and g665 (n_4771, n_4735, n_4375);
  or g666 (n_4775, n_4771, n_4772);
  and g667 (n_4773, n_4737, n_4375);
  or g668 (n_4776, n_4773, n_4774);
  and g669 (n_4778, n_4775, enT3);
  and g670 (n_4787, n_4776, enT3);
  and g671 (n_4802, n_4795, \Nanod[dbl2rxl] );
  and g672 (n_4799, n_4795, abdIsByte);
  and g673 (n_4798, n_4795, n_4318);
  or g674 (n_4800, n_4798, n_4799);
  and g676 (n_4801, n_4800, n_4322);
  or g677 (n_4805, n_4801, n_4802);
  and g678 (n_4804, n_4798, n_4322);
  or g679 (n_4806, n_4804, n_4802);
  and g680 (n_4809, n_4805, n_525);
  and g681 (n_4811, n_4806, n_525);
  and g682 (n_4808, n_4795, rxIsAreg);
  or g683 (n_4812, n_4808, n_4809);
  or g685 (n_4813, n_4808, n_4811);
  and g686 (n_4814, n_4812, n_524);
  and g687 (n_4816, n_4813, n_524);
  and g688 (n_4815, n_4814, n_900);
  or g689 (n_4818, n_4815, n_899);
  and g690 (n_4817, n_4816, n_900);
  or g691 (n_4819, n_4817, n_899);
  and g692 (n_4834, n_4818, \Nanod[dbl2ryl] );
  and g693 (n_4837, n_4819, \Nanod[dbl2ryl] );
  and g699 (n_4828, n_4818, abdIsByte);
  and g700 (n_4831, n_4816, abdIsByte);
  and g705 (n_4827, n_4818, n_4318);
  or g706 (n_4832, n_4827, n_4828);
  and g707 (n_4830, n_4819, n_4318);
  or g708 (n_4835, n_4830, n_4831);
  and g709 (n_4833, n_4832, n_4356);
  or g710 (n_4838, n_4833, n_4834);
  and g711 (n_4836, n_4835, n_4356);
  or g712 (n_4839, n_4836, n_4837);
  and g713 (n_4844, n_4838, n_521);
  and g714 (n_4847, n_4839, n_521);
  and g719 (n_4843, n_4818, ryIsAreg);
  or g720 (n_4848, n_4843, n_4844);
  and g721 (n_4846, n_4819, ryIsAreg);
  or g722 (n_4849, n_4846, n_4847);
  and g723 (n_4851, n_4848, n_520);
  and g724 (n_4853, n_4849, n_520);
  and g725 (n_4850, n_4814, n_4375);
  or g726 (n_4854, n_4850, n_4851);
  and g727 (n_4852, n_4816, n_4375);
  or g728 (n_4855, n_4852, n_4853);
  and g729 (n_4857, n_4854, enT3);
  and g730 (n_4866, n_4855, enT3);
  and g731 (n_4881, n_4874, \Nanod[dbl2rxl] );
  and g732 (n_4878, n_4874, abdIsByte);
  and g733 (n_4877, n_4874, n_4318);
  or g734 (n_4879, n_4877, n_4878);
  and g736 (n_4880, n_4879, n_4322);
  or g737 (n_4884, n_4880, n_4881);
  and g738 (n_4883, n_4877, n_4322);
  or g739 (n_4885, n_4883, n_4881);
  and g740 (n_4888, n_4884, n_525);
  and g741 (n_4890, n_4885, n_525);
  and g742 (n_4887, n_4874, rxIsAreg);
  or g743 (n_4891, n_4887, n_4888);
  or g745 (n_4892, n_4887, n_4890);
  and g746 (n_4893, n_4891, n_524);
  and g747 (n_4895, n_4892, n_524);
  and g748 (n_4894, n_4893, n_882);
  or g749 (n_4897, n_4894, n_881);
  and g750 (n_4896, n_4895, n_882);
  or g751 (n_4898, n_4896, n_881);
  and g752 (n_4913, n_4897, \Nanod[dbl2ryl] );
  and g753 (n_4916, n_4898, \Nanod[dbl2ryl] );
  and g759 (n_4907, n_4897, abdIsByte);
  and g760 (n_4910, n_4895, abdIsByte);
  and g765 (n_4906, n_4897, n_4318);
  or g766 (n_4911, n_4906, n_4907);
  and g767 (n_4909, n_4898, n_4318);
  or g768 (n_4914, n_4909, n_4910);
  and g769 (n_4912, n_4911, n_4356);
  or g770 (n_4917, n_4912, n_4913);
  and g771 (n_4915, n_4914, n_4356);
  or g772 (n_4918, n_4915, n_4916);
  and g773 (n_4923, n_4917, n_521);
  and g774 (n_4926, n_4918, n_521);
  and g779 (n_4922, n_4897, ryIsAreg);
  or g780 (n_4927, n_4922, n_4923);
  and g781 (n_4925, n_4898, ryIsAreg);
  or g782 (n_4928, n_4925, n_4926);
  and g783 (n_4930, n_4927, n_520);
  and g784 (n_4932, n_4928, n_520);
  and g785 (n_4929, n_4893, n_4375);
  or g786 (n_4933, n_4929, n_4930);
  and g787 (n_4931, n_4895, n_4375);
  or g788 (n_4934, n_4931, n_4932);
  and g789 (n_4936, n_4933, enT3);
  and g790 (n_4945, n_4934, enT3);
  and g791 (n_4960, n_4953, \Nanod[dbl2rxl] );
  and g792 (n_4957, n_4953, abdIsByte);
  and g793 (n_4956, n_4953, n_4318);
  or g794 (n_4958, n_4956, n_4957);
  and g796 (n_4959, n_4958, n_4322);
  or g797 (n_4963, n_4959, n_4960);
  and g798 (n_4962, n_4956, n_4322);
  or g799 (n_4964, n_4962, n_4960);
  and g800 (n_4967, n_4963, n_525);
  and g801 (n_4969, n_4964, n_525);
  and g802 (n_4966, n_4953, rxIsAreg);
  or g803 (n_4970, n_4966, n_4967);
  or g805 (n_4971, n_4966, n_4969);
  and g806 (n_4972, n_4970, n_524);
  and g807 (n_4974, n_4971, n_524);
  and g808 (n_4973, n_4972, n_864);
  or g809 (n_4976, n_4973, n_863);
  and g810 (n_4975, n_4974, n_864);
  or g811 (n_4977, n_4975, n_863);
  and g812 (n_4992, n_4976, \Nanod[dbl2ryl] );
  and g813 (n_4995, n_4977, \Nanod[dbl2ryl] );
  and g819 (n_4986, n_4976, abdIsByte);
  and g820 (n_4989, n_4974, abdIsByte);
  and g825 (n_4985, n_4976, n_4318);
  or g826 (n_4990, n_4985, n_4986);
  and g827 (n_4988, n_4977, n_4318);
  or g828 (n_4993, n_4988, n_4989);
  and g829 (n_4991, n_4990, n_4356);
  or g830 (n_4996, n_4991, n_4992);
  and g831 (n_4994, n_4993, n_4356);
  or g832 (n_4997, n_4994, n_4995);
  and g833 (n_5002, n_4996, n_521);
  and g834 (n_5005, n_4997, n_521);
  and g839 (n_5001, n_4976, ryIsAreg);
  or g840 (n_5006, n_5001, n_5002);
  and g841 (n_5004, n_4977, ryIsAreg);
  or g842 (n_5007, n_5004, n_5005);
  and g843 (n_5009, n_5006, n_520);
  and g844 (n_5011, n_5007, n_520);
  and g845 (n_5008, n_4972, n_4375);
  or g846 (n_5012, n_5008, n_5009);
  and g847 (n_5010, n_4974, n_4375);
  or g848 (n_5013, n_5010, n_5011);
  and g849 (n_5015, n_5012, enT3);
  and g850 (n_5024, n_5013, enT3);
  and g851 (n_5039, n_5032, \Nanod[dbl2rxl] );
  and g852 (n_5036, n_5032, abdIsByte);
  and g853 (n_5035, n_5032, n_4318);
  or g854 (n_5037, n_5035, n_5036);
  and g856 (n_5038, n_5037, n_4322);
  or g857 (n_5042, n_5038, n_5039);
  and g858 (n_5041, n_5035, n_4322);
  or g859 (n_5043, n_5041, n_5039);
  and g860 (n_5046, n_5042, n_525);
  and g861 (n_5048, n_5043, n_525);
  and g862 (n_5045, n_5032, rxIsAreg);
  or g863 (n_5049, n_5045, n_5046);
  or g865 (n_5050, n_5045, n_5048);
  and g866 (n_5051, n_5049, n_524);
  and g867 (n_5053, n_5050, n_524);
  and g868 (n_5052, n_5051, n_846);
  or g869 (n_5055, n_5052, n_845);
  and g870 (n_5054, n_5053, n_846);
  or g871 (n_5056, n_5054, n_845);
  and g872 (n_5071, n_5055, \Nanod[dbl2ryl] );
  and g873 (n_5074, n_5056, \Nanod[dbl2ryl] );
  and g879 (n_5065, n_5055, abdIsByte);
  and g880 (n_5068, n_5053, abdIsByte);
  and g885 (n_5064, n_5055, n_4318);
  or g886 (n_5069, n_5064, n_5065);
  and g887 (n_5067, n_5056, n_4318);
  or g888 (n_5072, n_5067, n_5068);
  and g889 (n_5070, n_5069, n_4356);
  or g890 (n_5075, n_5070, n_5071);
  and g891 (n_5073, n_5072, n_4356);
  or g892 (n_5076, n_5073, n_5074);
  and g893 (n_5081, n_5075, n_521);
  and g894 (n_5084, n_5076, n_521);
  and g899 (n_5080, n_5055, ryIsAreg);
  or g900 (n_5085, n_5080, n_5081);
  and g901 (n_5083, n_5056, ryIsAreg);
  or g902 (n_5086, n_5083, n_5084);
  and g903 (n_5088, n_5085, n_520);
  and g904 (n_5090, n_5086, n_520);
  and g905 (n_5087, n_5051, n_4375);
  or g906 (n_5091, n_5087, n_5088);
  and g907 (n_5089, n_5053, n_4375);
  or g908 (n_5092, n_5089, n_5090);
  and g909 (n_5094, n_5091, enT3);
  and g910 (n_5103, n_5092, enT3);
  and g911 (n_5118, n_5111, \Nanod[dbl2rxl] );
  and g912 (n_5115, n_5111, abdIsByte);
  and g913 (n_5114, n_5111, n_4318);
  or g914 (n_5116, n_5114, n_5115);
  and g916 (n_5117, n_5116, n_4322);
  or g917 (n_5121, n_5117, n_5118);
  and g918 (n_5120, n_5114, n_4322);
  or g919 (n_5122, n_5120, n_5118);
  and g920 (n_5125, n_5121, n_525);
  and g921 (n_5127, n_5122, n_525);
  and g922 (n_5124, n_5111, rxIsAreg);
  or g923 (n_5128, n_5124, n_5125);
  or g925 (n_5129, n_5124, n_5127);
  and g926 (n_5130, n_5128, n_524);
  and g927 (n_5132, n_5129, n_524);
  and g928 (n_5131, n_5130, n_828);
  or g929 (n_5134, n_5131, n_827);
  and g930 (n_5133, n_5132, n_828);
  or g931 (n_5135, n_5133, n_827);
  and g932 (n_5150, n_5134, \Nanod[dbl2ryl] );
  and g933 (n_5153, n_5135, \Nanod[dbl2ryl] );
  and g939 (n_5144, n_5134, abdIsByte);
  and g940 (n_5147, n_5132, abdIsByte);
  and g945 (n_5143, n_5134, n_4318);
  or g946 (n_5148, n_5143, n_5144);
  and g947 (n_5146, n_5135, n_4318);
  or g948 (n_5151, n_5146, n_5147);
  and g949 (n_5149, n_5148, n_4356);
  or g950 (n_5154, n_5149, n_5150);
  and g951 (n_5152, n_5151, n_4356);
  or g952 (n_5155, n_5152, n_5153);
  and g953 (n_5160, n_5154, n_521);
  and g954 (n_5163, n_5155, n_521);
  and g959 (n_5159, n_5134, ryIsAreg);
  or g960 (n_5164, n_5159, n_5160);
  and g961 (n_5162, n_5135, ryIsAreg);
  or g962 (n_5165, n_5162, n_5163);
  and g963 (n_5167, n_5164, n_520);
  and g964 (n_5169, n_5165, n_520);
  and g965 (n_5166, n_5130, n_4375);
  or g966 (n_5170, n_5166, n_5167);
  and g967 (n_5168, n_5132, n_4375);
  or g968 (n_5171, n_5168, n_5169);
  and g969 (n_5173, n_5170, enT3);
  and g970 (n_5182, n_5171, enT3);
  and g971 (n_5197, n_5190, \Nanod[dbl2rxl] );
  and g972 (n_5194, n_5190, abdIsByte);
  and g973 (n_5193, n_5190, n_4318);
  or g974 (n_5195, n_5193, n_5194);
  and g976 (n_5196, n_5195, n_4322);
  or g977 (n_5200, n_5196, n_5197);
  and g978 (n_5199, n_5193, n_4322);
  or g979 (n_5201, n_5199, n_5197);
  and g980 (n_5204, n_5200, n_525);
  and g981 (n_5206, n_5201, n_525);
  and g982 (n_5203, n_5190, rxIsAreg);
  or g983 (n_5207, n_5203, n_5204);
  or g985 (n_5208, n_5203, n_5206);
  and g986 (n_5209, n_5207, n_524);
  and g987 (n_5211, n_5208, n_524);
  and g988 (n_5210, n_5209, n_810);
  or g989 (n_5213, n_5210, n_809);
  and g990 (n_5212, n_5211, n_810);
  or g991 (n_5214, n_5212, n_809);
  and g992 (n_5229, n_5213, \Nanod[dbl2ryl] );
  and g993 (n_5232, n_5214, \Nanod[dbl2ryl] );
  and g999 (n_5223, n_5213, abdIsByte);
  and g1000 (n_5226, n_5211, abdIsByte);
  and g1005 (n_5222, n_5213, n_4318);
  or g1006 (n_5227, n_5222, n_5223);
  and g1007 (n_5225, n_5214, n_4318);
  or g1008 (n_5230, n_5225, n_5226);
  and g1009 (n_5228, n_5227, n_4356);
  or g1010 (n_5233, n_5228, n_5229);
  and g1011 (n_5231, n_5230, n_4356);
  or g1012 (n_5234, n_5231, n_5232);
  and g1013 (n_5239, n_5233, n_521);
  and g1014 (n_5242, n_5234, n_521);
  and g1019 (n_5238, n_5213, ryIsAreg);
  or g1020 (n_5243, n_5238, n_5239);
  and g1021 (n_5241, n_5214, ryIsAreg);
  or g1022 (n_5244, n_5241, n_5242);
  and g1023 (n_5246, n_5243, n_520);
  and g1024 (n_5248, n_5244, n_520);
  and g1025 (n_5245, n_5209, n_4375);
  or g1026 (n_5249, n_5245, n_5246);
  and g1027 (n_5247, n_5211, n_4375);
  or g1028 (n_5250, n_5247, n_5248);
  and g1029 (n_5252, n_5249, enT3);
  and g1030 (n_5261, n_5250, enT3);
  and g1031 (n_5276, n_5269, \Nanod[dbl2rxl] );
  and g1032 (n_5273, n_5269, abdIsByte);
  and g1033 (n_5272, n_5269, n_4318);
  or g1034 (n_5274, n_5272, n_5273);
  and g1036 (n_5275, n_5274, n_4322);
  or g1037 (n_5279, n_5275, n_5276);
  and g1038 (n_5278, n_5272, n_4322);
  or g1039 (n_5280, n_5278, n_5276);
  and g1040 (n_5283, n_5279, n_525);
  and g1041 (n_5285, n_5280, n_525);
  and g1042 (n_5282, n_5269, rxIsAreg);
  or g1043 (n_5286, n_5282, n_5283);
  or g1045 (n_5287, n_5282, n_5285);
  and g1046 (n_5288, n_5286, n_524);
  and g1047 (n_5290, n_5287, n_524);
  and g1048 (n_5289, n_5288, n_792);
  or g1049 (n_5292, n_5289, n_791);
  and g1050 (n_5291, n_5290, n_792);
  or g1051 (n_5293, n_5291, n_791);
  and g1052 (n_5308, n_5292, \Nanod[dbl2ryl] );
  and g1053 (n_5311, n_5293, \Nanod[dbl2ryl] );
  and g1059 (n_5302, n_5292, abdIsByte);
  and g1060 (n_5305, n_5290, abdIsByte);
  and g1065 (n_5301, n_5292, n_4318);
  or g1066 (n_5306, n_5301, n_5302);
  and g1067 (n_5304, n_5293, n_4318);
  or g1068 (n_5309, n_5304, n_5305);
  and g1069 (n_5307, n_5306, n_4356);
  or g1070 (n_5312, n_5307, n_5308);
  and g1071 (n_5310, n_5309, n_4356);
  or g1072 (n_5313, n_5310, n_5311);
  and g1073 (n_5318, n_5312, n_521);
  and g1074 (n_5321, n_5313, n_521);
  and g1079 (n_5317, n_5292, ryIsAreg);
  or g1080 (n_5322, n_5317, n_5318);
  and g1081 (n_5320, n_5293, ryIsAreg);
  or g1082 (n_5323, n_5320, n_5321);
  and g1083 (n_5325, n_5322, n_520);
  and g1084 (n_5327, n_5323, n_520);
  and g1085 (n_5324, n_5288, n_4375);
  or g1086 (n_5328, n_5324, n_5325);
  and g1087 (n_5326, n_5290, n_4375);
  or g1088 (n_5329, n_5326, n_5327);
  and g1089 (n_5331, n_5328, enT3);
  and g1090 (n_5340, n_5329, enT3);
  and g1091 (n_5355, n_5348, \Nanod[dbl2rxl] );
  and g1092 (n_5352, n_5348, abdIsByte);
  and g1093 (n_5351, n_5348, n_4318);
  or g1094 (n_5353, n_5351, n_5352);
  and g1096 (n_5354, n_5353, n_4322);
  or g1097 (n_5358, n_5354, n_5355);
  and g1098 (n_5357, n_5351, n_4322);
  or g1099 (n_5359, n_5357, n_5355);
  and g1100 (n_5362, n_5358, n_525);
  and g1101 (n_5364, n_5359, n_525);
  and g1102 (n_5361, n_5348, rxIsAreg);
  or g1103 (n_5365, n_5361, n_5362);
  or g1105 (n_5366, n_5361, n_5364);
  and g1106 (n_5367, n_5365, n_524);
  and g1107 (n_5369, n_5366, n_524);
  and g1108 (n_5368, n_5367, n_774);
  or g1109 (n_5371, n_5368, n_773);
  and g1110 (n_5370, n_5369, n_774);
  or g1111 (n_5372, n_5370, n_773);
  and g1112 (n_5387, n_5371, \Nanod[dbl2ryl] );
  and g1113 (n_5390, n_5372, \Nanod[dbl2ryl] );
  and g1119 (n_5381, n_5371, abdIsByte);
  and g1120 (n_5384, n_5369, abdIsByte);
  and g1125 (n_5380, n_5371, n_4318);
  or g1126 (n_5385, n_5380, n_5381);
  and g1127 (n_5383, n_5372, n_4318);
  or g1128 (n_5388, n_5383, n_5384);
  and g1129 (n_5386, n_5385, n_4356);
  or g1130 (n_5391, n_5386, n_5387);
  and g1131 (n_5389, n_5388, n_4356);
  or g1132 (n_5392, n_5389, n_5390);
  and g1133 (n_5397, n_5391, n_521);
  and g1134 (n_5400, n_5392, n_521);
  and g1139 (n_5396, n_5371, ryIsAreg);
  or g1140 (n_5401, n_5396, n_5397);
  and g1141 (n_5399, n_5372, ryIsAreg);
  or g1142 (n_5402, n_5399, n_5400);
  and g1143 (n_5404, n_5401, n_520);
  and g1144 (n_5406, n_5402, n_520);
  and g1145 (n_5403, n_5367, n_4375);
  or g1146 (n_5407, n_5403, n_5404);
  and g1147 (n_5405, n_5369, n_4375);
  or g1148 (n_5408, n_5405, n_5406);
  and g1149 (n_5410, n_5407, enT3);
  and g1150 (n_5419, n_5408, enT3);
  and g1151 (n_5434, n_5427, \Nanod[dbl2rxl] );
  and g1152 (n_5431, n_5427, abdIsByte);
  and g1153 (n_5430, n_5427, n_4318);
  or g1154 (n_5432, n_5430, n_5431);
  and g1156 (n_5433, n_5432, n_4322);
  or g1157 (n_5437, n_5433, n_5434);
  and g1158 (n_5436, n_5430, n_4322);
  or g1159 (n_5438, n_5436, n_5434);
  and g1160 (n_5441, n_5437, n_525);
  and g1161 (n_5443, n_5438, n_525);
  and g1162 (n_5440, n_5427, rxIsAreg);
  or g1163 (n_5444, n_5440, n_5441);
  or g1165 (n_5445, n_5440, n_5443);
  and g1166 (n_5446, n_5444, n_524);
  and g1167 (n_5448, n_5445, n_524);
  and g1168 (n_5447, n_5446, n_756);
  or g1169 (n_5450, n_5447, n_755);
  and g1170 (n_5449, n_5448, n_756);
  or g1171 (n_5451, n_5449, n_755);
  and g1172 (n_5466, n_5450, \Nanod[dbl2ryl] );
  and g1173 (n_5469, n_5451, \Nanod[dbl2ryl] );
  and g1179 (n_5460, n_5450, abdIsByte);
  and g1180 (n_5463, n_5448, abdIsByte);
  and g1185 (n_5459, n_5450, n_4318);
  or g1186 (n_5464, n_5459, n_5460);
  and g1187 (n_5462, n_5451, n_4318);
  or g1188 (n_5467, n_5462, n_5463);
  and g1189 (n_5465, n_5464, n_4356);
  or g1190 (n_5470, n_5465, n_5466);
  and g1191 (n_5468, n_5467, n_4356);
  or g1192 (n_5471, n_5468, n_5469);
  and g1193 (n_5476, n_5470, n_521);
  and g1194 (n_5479, n_5471, n_521);
  and g1199 (n_5475, n_5450, ryIsAreg);
  or g1200 (n_5480, n_5475, n_5476);
  and g1201 (n_5478, n_5451, ryIsAreg);
  or g1202 (n_5481, n_5478, n_5479);
  and g1203 (n_5483, n_5480, n_520);
  and g1204 (n_5485, n_5481, n_520);
  and g1205 (n_5482, n_5446, n_4375);
  or g1206 (n_5486, n_5482, n_5483);
  and g1207 (n_5484, n_5448, n_4375);
  or g1208 (n_5487, n_5484, n_5485);
  and g1209 (n_5489, n_5486, enT3);
  and g1210 (n_5498, n_5487, enT3);
  and g1211 (n_5513, n_5506, \Nanod[dbl2rxl] );
  and g1212 (n_5510, n_5506, abdIsByte);
  and g1213 (n_5509, n_5506, n_4318);
  or g1214 (n_5511, n_5509, n_5510);
  and g1216 (n_5512, n_5511, n_4322);
  or g1217 (n_5516, n_5512, n_5513);
  and g1218 (n_5515, n_5509, n_4322);
  or g1219 (n_5517, n_5515, n_5513);
  and g1220 (n_5520, n_5516, n_525);
  and g1221 (n_5522, n_5517, n_525);
  and g1222 (n_5519, n_5506, rxIsAreg);
  or g1223 (n_5523, n_5519, n_5520);
  or g1225 (n_5524, n_5519, n_5522);
  and g1226 (n_5525, n_5523, n_524);
  and g1227 (n_5527, n_5524, n_524);
  and g1228 (n_5526, n_5525, n_738);
  or g1229 (n_5529, n_5526, n_737);
  and g1230 (n_5528, n_5527, n_738);
  or g1231 (n_5530, n_5528, n_737);
  and g1232 (n_5545, n_5529, \Nanod[dbl2ryl] );
  and g1233 (n_5548, n_5530, \Nanod[dbl2ryl] );
  and g1239 (n_5539, n_5529, abdIsByte);
  and g1240 (n_5542, n_5527, abdIsByte);
  and g1245 (n_5538, n_5529, n_4318);
  or g1246 (n_5543, n_5538, n_5539);
  and g1247 (n_5541, n_5530, n_4318);
  or g1248 (n_5546, n_5541, n_5542);
  and g1249 (n_5544, n_5543, n_4356);
  or g1250 (n_5549, n_5544, n_5545);
  and g1251 (n_5547, n_5546, n_4356);
  or g1252 (n_5550, n_5547, n_5548);
  and g1253 (n_5555, n_5549, n_521);
  and g1254 (n_5558, n_5550, n_521);
  and g1259 (n_5554, n_5529, ryIsAreg);
  or g1260 (n_5559, n_5554, n_5555);
  and g1261 (n_5557, n_5530, ryIsAreg);
  or g1262 (n_5560, n_5557, n_5558);
  and g1263 (n_5562, n_5559, n_520);
  and g1264 (n_5564, n_5560, n_520);
  and g1265 (n_5561, n_5525, n_4375);
  or g1266 (n_5565, n_5561, n_5562);
  and g1267 (n_5563, n_5527, n_4375);
  or g1268 (n_5566, n_5563, n_5564);
  and g1269 (n_5568, n_5565, enT3);
  and g1270 (n_5577, n_5566, enT3);
  and g1271 (n_5592, n_5585, \Nanod[dbl2rxl] );
  and g1272 (n_5589, n_5585, abdIsByte);
  and g1273 (n_5588, n_5585, n_4318);
  or g1274 (n_5590, n_5588, n_5589);
  and g1276 (n_5591, n_5590, n_4322);
  or g1277 (n_5595, n_5591, n_5592);
  and g1278 (n_5594, n_5588, n_4322);
  or g1279 (n_5596, n_5594, n_5592);
  and g1280 (n_5599, n_5595, n_525);
  and g1281 (n_5601, n_5596, n_525);
  and g1282 (n_5598, n_5585, rxIsAreg);
  or g1283 (n_5602, n_5598, n_5599);
  or g1285 (n_5603, n_5598, n_5601);
  and g1286 (n_5604, n_5602, n_524);
  and g1287 (n_5606, n_5603, n_524);
  and g1288 (n_5605, n_5604, n_720);
  or g1289 (n_5608, n_5605, n_719);
  and g1290 (n_5607, n_5606, n_720);
  or g1291 (n_5609, n_5607, n_719);
  and g1292 (n_5624, n_5608, \Nanod[dbl2ryl] );
  and g1293 (n_5627, n_5609, \Nanod[dbl2ryl] );
  and g1299 (n_5618, n_5608, abdIsByte);
  and g1300 (n_5621, n_5606, abdIsByte);
  and g1305 (n_5617, n_5608, n_4318);
  or g1306 (n_5622, n_5617, n_5618);
  and g1307 (n_5620, n_5609, n_4318);
  or g1308 (n_5625, n_5620, n_5621);
  and g1309 (n_5623, n_5622, n_4356);
  or g1310 (n_5628, n_5623, n_5624);
  and g1311 (n_5626, n_5625, n_4356);
  or g1312 (n_5629, n_5626, n_5627);
  and g1313 (n_5634, n_5628, n_521);
  and g1314 (n_5637, n_5629, n_521);
  and g1319 (n_5633, n_5608, ryIsAreg);
  or g1320 (n_5638, n_5633, n_5634);
  and g1321 (n_5636, n_5609, ryIsAreg);
  or g1322 (n_5639, n_5636, n_5637);
  and g1323 (n_5641, n_5638, n_520);
  and g1324 (n_5643, n_5639, n_520);
  and g1325 (n_5640, n_5604, n_4375);
  or g1326 (n_5644, n_5640, n_5641);
  and g1327 (n_5642, n_5606, n_4375);
  or g1328 (n_5645, n_5642, n_5643);
  and g1329 (n_5647, n_5644, enT3);
  and g1330 (n_5656, n_5645, enT3);
  and g1331 (n_5671, n_5664, \Nanod[dbl2rxl] );
  and g1332 (n_5668, n_5664, abdIsByte);
  and g1333 (n_5667, n_5664, n_4318);
  or g1334 (n_5669, n_5667, n_5668);
  and g1336 (n_5670, n_5669, n_4322);
  or g1337 (n_5674, n_5670, n_5671);
  and g1338 (n_5673, n_5667, n_4322);
  or g1339 (n_5675, n_5673, n_5671);
  and g1340 (n_5678, n_5674, n_525);
  and g1341 (n_5680, n_5675, n_525);
  and g1342 (n_5677, n_5664, rxIsAreg);
  or g1343 (n_5681, n_5677, n_5678);
  or g1345 (n_5682, n_5677, n_5680);
  and g1346 (n_5683, n_5681, n_524);
  and g1347 (n_5685, n_5682, n_524);
  and g1348 (n_5684, n_5683, n_670);
  or g1349 (n_5687, n_5684, n_669);
  and g1350 (n_5686, n_5685, n_670);
  or g1351 (n_5688, n_5686, n_669);
  and g1352 (n_5703, n_5687, \Nanod[dbl2ryl] );
  and g1353 (n_5706, n_5688, \Nanod[dbl2ryl] );
  and g1359 (n_5697, n_5687, abdIsByte);
  and g1360 (n_5700, n_5685, abdIsByte);
  and g1365 (n_5696, n_5687, n_4318);
  or g1366 (n_5701, n_5696, n_5697);
  and g1367 (n_5699, n_5688, n_4318);
  or g1368 (n_5704, n_5699, n_5700);
  and g1369 (n_5702, n_5701, n_4356);
  or g1370 (n_5707, n_5702, n_5703);
  and g1371 (n_5705, n_5704, n_4356);
  or g1372 (n_5708, n_5705, n_5706);
  and g1373 (n_5713, n_5707, n_521);
  and g1374 (n_5716, n_5708, n_521);
  and g1379 (n_5712, n_5687, ryIsAreg);
  or g1380 (n_5717, n_5712, n_5713);
  and g1381 (n_5715, n_5688, ryIsAreg);
  or g1382 (n_5718, n_5715, n_5716);
  and g1383 (n_5720, n_5717, n_520);
  and g1384 (n_5722, n_5718, n_520);
  and g1385 (n_5719, n_5683, n_4375);
  or g1386 (n_5723, n_5719, n_5720);
  and g1387 (n_5721, n_5685, n_4375);
  or g1388 (n_5724, n_5721, n_5722);
  and g1389 (n_5726, n_5723, enT3);
  and g1390 (n_5735, n_5724, enT3);
  and g1391 (n_5744, n_4315, n_667);
  and g1392 (n_5745, n_5744, n_1008);
  or g1393 (n_5746, n_5745, n_1007);
  and g1394 (n_5749, n_5746, n_654);
  and g1395 (n_5748, n_5744, n_5747);
  or g1396 (n_5750, n_5748, n_5749);
  and g1397 (n_5752, n_5750, enT3);
  and g1398 (n_5769, n_4400, n_667);
  and g1399 (n_5770, n_5769, n_990);
  or g1400 (n_5771, n_5770, n_989);
  and g1401 (n_5773, n_5771, n_654);
  and g1402 (n_5772, n_5769, n_5747);
  or g1403 (n_5774, n_5772, n_5773);
  and g1404 (n_5776, n_5774, enT3);
  and g1405 (n_5793, n_4479, n_667);
  and g1406 (n_5794, n_5793, n_972);
  or g1407 (n_5795, n_5794, n_971);
  and g1408 (n_5797, n_5795, n_654);
  and g1409 (n_5796, n_5793, n_5747);
  or g1410 (n_5798, n_5796, n_5797);
  and g1411 (n_5800, n_5798, enT3);
  and g1412 (n_5817, n_4558, n_667);
  and g1413 (n_5818, n_5817, n_954);
  or g1414 (n_5819, n_5818, n_953);
  and g1415 (n_5821, n_5819, n_654);
  and g1416 (n_5820, n_5817, n_5747);
  or g1417 (n_5822, n_5820, n_5821);
  and g1418 (n_5824, n_5822, enT3);
  and g1419 (n_5841, n_4637, n_667);
  and g1420 (n_5842, n_5841, n_936);
  or g1421 (n_5843, n_5842, n_935);
  and g1422 (n_5845, n_5843, n_654);
  and g1423 (n_5844, n_5841, n_5747);
  or g1424 (n_5846, n_5844, n_5845);
  and g1425 (n_5848, n_5846, enT3);
  and g1426 (n_5865, n_4716, n_667);
  and g1427 (n_5866, n_5865, n_918);
  or g1428 (n_5867, n_5866, n_917);
  and g1429 (n_5869, n_5867, n_654);
  and g1430 (n_5868, n_5865, n_5747);
  or g1431 (n_5870, n_5868, n_5869);
  and g1432 (n_5872, n_5870, enT3);
  and g1433 (n_5889, n_4795, n_667);
  and g1434 (n_5890, n_5889, n_900);
  or g1435 (n_5891, n_5890, n_899);
  and g1436 (n_5893, n_5891, n_654);
  and g1437 (n_5892, n_5889, n_5747);
  or g1438 (n_5894, n_5892, n_5893);
  and g1439 (n_5896, n_5894, enT3);
  and g1440 (n_5913, n_4874, n_667);
  and g1441 (n_5914, n_5913, n_882);
  or g1442 (n_5915, n_5914, n_881);
  and g1443 (n_5917, n_5915, n_654);
  and g1444 (n_5916, n_5913, n_5747);
  or g1445 (n_5918, n_5916, n_5917);
  and g1446 (n_5920, n_5918, enT3);
  and g1447 (n_5937, n_4953, n_667);
  and g1448 (n_5938, n_5937, n_864);
  or g1449 (n_5939, n_5938, n_863);
  and g1450 (n_5941, n_5939, n_654);
  and g1451 (n_5940, n_5937, n_5747);
  or g1452 (n_5942, n_5940, n_5941);
  and g1453 (n_5944, n_5942, enT3);
  and g1454 (n_5961, n_5032, n_667);
  and g1455 (n_5962, n_5961, n_846);
  or g1456 (n_5963, n_5962, n_845);
  and g1457 (n_5965, n_5963, n_654);
  and g1458 (n_5964, n_5961, n_5747);
  or g1459 (n_5966, n_5964, n_5965);
  and g1460 (n_5968, n_5966, enT3);
  and g1461 (n_5985, n_5111, n_667);
  and g1462 (n_5986, n_5985, n_828);
  or g1463 (n_5987, n_5986, n_827);
  and g1464 (n_5989, n_5987, n_654);
  and g1465 (n_5988, n_5985, n_5747);
  or g1466 (n_5990, n_5988, n_5989);
  and g1467 (n_5992, n_5990, enT3);
  and g1468 (n_6009, n_5190, n_667);
  and g1469 (n_6010, n_6009, n_810);
  or g1470 (n_6011, n_6010, n_809);
  and g1471 (n_6013, n_6011, n_654);
  and g1472 (n_6012, n_6009, n_5747);
  or g1473 (n_6014, n_6012, n_6013);
  and g1474 (n_6016, n_6014, enT3);
  and g1475 (n_6033, n_5269, n_667);
  and g1476 (n_6034, n_6033, n_792);
  or g1477 (n_6035, n_6034, n_791);
  and g1478 (n_6037, n_6035, n_654);
  and g1479 (n_6036, n_6033, n_5747);
  or g1480 (n_6038, n_6036, n_6037);
  and g1481 (n_6040, n_6038, enT3);
  and g1482 (n_6057, n_5348, n_667);
  and g1483 (n_6058, n_6057, n_774);
  or g1484 (n_6059, n_6058, n_773);
  and g1485 (n_6061, n_6059, n_654);
  and g1486 (n_6060, n_6057, n_5747);
  or g1487 (n_6062, n_6060, n_6061);
  and g1488 (n_6064, n_6062, enT3);
  and g1489 (n_6081, n_5427, n_667);
  and g1490 (n_6082, n_6081, n_756);
  or g1491 (n_6083, n_6082, n_755);
  and g1492 (n_6085, n_6083, n_654);
  and g1493 (n_6084, n_6081, n_5747);
  or g1494 (n_6086, n_6084, n_6085);
  and g1495 (n_6088, n_6086, enT3);
  and g1496 (n_6105, n_5506, n_667);
  and g1497 (n_6106, n_6105, n_738);
  or g1498 (n_6107, n_6106, n_737);
  and g1499 (n_6109, n_6107, n_654);
  and g1500 (n_6108, n_6105, n_5747);
  or g1501 (n_6110, n_6108, n_6109);
  and g1502 (n_6112, n_6110, enT3);
  and g1503 (n_6129, n_5585, n_667);
  and g1504 (n_6130, n_6129, n_720);
  or g1505 (n_6131, n_6130, n_719);
  and g1506 (n_6133, n_6131, n_654);
  and g1507 (n_6132, n_6129, n_5747);
  or g1508 (n_6134, n_6132, n_6133);
  and g1509 (n_6136, n_6134, enT3);
  and g1510 (n_6153, n_5664, n_667);
  and g1511 (n_6154, n_6153, n_670);
  or g1512 (n_6155, n_6154, n_669);
  and g1513 (n_6157, n_6155, n_654);
  and g1514 (n_6156, n_6153, n_5747);
  or g1515 (n_6158, n_6156, n_6157);
  and g1516 (n_6160, n_6158, enT3);
  and g1517 (n_6177, abl2Pcl, n_6176);
  or g1518 (n_6178, n_6177, dbl2Pcl);
  and g1519 (n_6179, n_6178, enT3);
  and g1520 (n_6181, n_6179, n_6180);
  or g1521 (n_6183, n_6181, n_553);
  and g1522 (n_6200, abh2Pch, n_6199);
  or g1523 (n_6201, n_6200, dbh2Pch);
  and g1524 (n_6202, n_6201, enT3);
  and g1525 (n_6204, n_6202, n_6180);
  or g1526 (n_6206, n_6204, n_553);
  and g1527 (n_6223, \Nanod[dbh2Ath] , n_6222);
  or g1528 (n_6224, n_6223, \Nanod[abh2Ath] );
  and g1529 (n_6226, n_6224, enT3);
  and g1530 (n_6243, \Nanod[abl2Atl] , n_6242);
  or g1531 (n_6244, n_6243, \Nanod[dbl2Atl] );
  and g1532 (n_6246, n_6244, enT3);
  and g1533 (n_6264, n_457, n_6262);
  or g1535 (n_6270, n_6264, n_456);
  and g1536 (n_6287, n_643, n_6286);
  and g1537 (n_6289, \Nanod[abd2Alub] , n_6288);
  or g1538 (n_6290, n_6289, \Nanod[dbd2Alub] );
  and g1539 (n_6292, n_6290, enT3);
  nor g1 (n_6351, auReg[5], auReg[4], auReg[3], auReg[2]);
  nor g1540 (n_6350, auReg[1], auReg[0]);
  nand g1541 (n_6352, n_6350, n_6351);
  not g1542 (au05z, n_6352);
  not g1543 (n_4178, \Irdecod[implicitSp] );
  not g1544 (n_4179, \Nanod[rz] );
  CDN_flop abdIsByte_reg(.clk (\Clks[clk] ), .d (n_4183), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (abdIsByte));
  CDN_flop \actualRx_reg[0] (.clk (\Clks[clk] ), .d (rxMux[0]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRx[0]));
  CDN_flop \actualRx_reg[1] (.clk (\Clks[clk] ), .d (rxMux[1]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRx[1]));
  CDN_flop \actualRx_reg[2] (.clk (\Clks[clk] ), .d (rxMux[2]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRx[2]));
  CDN_flop \actualRx_reg[3] (.clk (\Clks[clk] ), .d (rxMux[3]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRx[3]));
  CDN_flop \actualRx_reg[4] (.clk (\Clks[clk] ), .d (rxMux[4]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRx[4]));
  CDN_flop \actualRy_reg[0] (.clk (\Clks[clk] ), .d (ryMux[0]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRy[0]));
  CDN_flop \actualRy_reg[1] (.clk (\Clks[clk] ), .d (ryMux[1]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRy[1]));
  CDN_flop \actualRy_reg[2] (.clk (\Clks[clk] ), .d (ryMux[2]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRy[2]));
  CDN_flop \actualRy_reg[3] (.clk (\Clks[clk] ), .d (ryMux[3]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRy[3]));
  CDN_flop \actualRy_reg[4] (.clk (\Clks[clk] ), .d (ryMux[4]), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (actualRy[4]));
  CDN_flop byteNotSpAlign_reg(.clk (\Clks[clk] ), .d (n_4184), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (byteNotSpAlign));
  CDN_flop rxIsAreg_reg(.clk (\Clks[clk] ), .d (n_4185), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (rxIsAreg));
  CDN_flop ryIsAreg_reg(.clk (\Clks[clk] ), .d (n_4186), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ryIsAreg));
  CDN_flop \Dbl_reg[0] (.clk (\Clks[clk] ), .d (n_4195), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[0]));
  CDN_flop \Dbl_reg[1] (.clk (\Clks[clk] ), .d (n_4196), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[1]));
  CDN_flop \Dbl_reg[2] (.clk (\Clks[clk] ), .d (n_4197), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[2]));
  CDN_flop \Dbl_reg[3] (.clk (\Clks[clk] ), .d (n_4198), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[3]));
  CDN_flop \Dbl_reg[4] (.clk (\Clks[clk] ), .d (n_4199), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[4]));
  CDN_flop \Dbl_reg[5] (.clk (\Clks[clk] ), .d (n_4200), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[5]));
  CDN_flop \Dbl_reg[6] (.clk (\Clks[clk] ), .d (n_4201), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[6]));
  CDN_flop \Dbl_reg[7] (.clk (\Clks[clk] ), .d (n_4202), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[7]));
  CDN_flop \Dbl_reg[8] (.clk (\Clks[clk] ), .d (n_4203), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[8]));
  CDN_flop \Dbl_reg[9] (.clk (\Clks[clk] ), .d (n_4204), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[9]));
  CDN_flop \Dbl_reg[10] (.clk (\Clks[clk] ), .d (n_4205), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[10]));
  CDN_flop \Dbl_reg[11] (.clk (\Clks[clk] ), .d (n_4206), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[11]));
  CDN_flop \Dbl_reg[12] (.clk (\Clks[clk] ), .d (n_4207), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[12]));
  CDN_flop \Dbl_reg[13] (.clk (\Clks[clk] ), .d (n_4208), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[13]));
  CDN_flop \Dbl_reg[14] (.clk (\Clks[clk] ), .d (n_4209), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[14]));
  CDN_flop \Dbl_reg[15] (.clk (\Clks[clk] ), .d (n_4210), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbl[15]));
  CDN_flop \Dbh_reg[0] (.clk (\Clks[clk] ), .d (n_4211), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[0]));
  CDN_flop \Dbh_reg[1] (.clk (\Clks[clk] ), .d (n_4212), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[1]));
  CDN_flop \Dbh_reg[2] (.clk (\Clks[clk] ), .d (n_4213), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[2]));
  CDN_flop \Dbh_reg[3] (.clk (\Clks[clk] ), .d (n_4214), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[3]));
  CDN_flop \Dbh_reg[4] (.clk (\Clks[clk] ), .d (n_4215), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[4]));
  CDN_flop \Dbh_reg[5] (.clk (\Clks[clk] ), .d (n_4216), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[5]));
  CDN_flop \Dbh_reg[6] (.clk (\Clks[clk] ), .d (n_4217), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[6]));
  CDN_flop \Dbh_reg[7] (.clk (\Clks[clk] ), .d (n_4218), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[7]));
  CDN_flop \Dbh_reg[8] (.clk (\Clks[clk] ), .d (n_4219), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[8]));
  CDN_flop \Dbh_reg[9] (.clk (\Clks[clk] ), .d (n_4220), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[9]));
  CDN_flop \Dbh_reg[10] (.clk (\Clks[clk] ), .d (n_4221), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[10]));
  CDN_flop \Dbh_reg[11] (.clk (\Clks[clk] ), .d (n_4222), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[11]));
  CDN_flop \Dbh_reg[12] (.clk (\Clks[clk] ), .d (n_4223), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[12]));
  CDN_flop \Dbh_reg[13] (.clk (\Clks[clk] ), .d (n_4224), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[13]));
  CDN_flop \Dbh_reg[14] (.clk (\Clks[clk] ), .d (n_4225), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[14]));
  CDN_flop \Dbh_reg[15] (.clk (\Clks[clk] ), .d (n_4226), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbh[15]));
  CDN_flop \Abh_reg[0] (.clk (\Clks[clk] ), .d (n_4227), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[0]));
  CDN_flop \Abh_reg[1] (.clk (\Clks[clk] ), .d (n_4228), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[1]));
  CDN_flop \Abh_reg[2] (.clk (\Clks[clk] ), .d (n_4229), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[2]));
  CDN_flop \Abh_reg[3] (.clk (\Clks[clk] ), .d (n_4230), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[3]));
  CDN_flop \Abh_reg[4] (.clk (\Clks[clk] ), .d (n_4231), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[4]));
  CDN_flop \Abh_reg[5] (.clk (\Clks[clk] ), .d (n_4232), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[5]));
  CDN_flop \Abh_reg[6] (.clk (\Clks[clk] ), .d (n_4233), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[6]));
  CDN_flop \Abh_reg[7] (.clk (\Clks[clk] ), .d (n_4234), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[7]));
  CDN_flop \Abh_reg[8] (.clk (\Clks[clk] ), .d (n_4235), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[8]));
  CDN_flop \Abh_reg[9] (.clk (\Clks[clk] ), .d (n_4236), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[9]));
  CDN_flop \Abh_reg[10] (.clk (\Clks[clk] ), .d (n_4237), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[10]));
  CDN_flop \Abh_reg[11] (.clk (\Clks[clk] ), .d (n_4238), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[11]));
  CDN_flop \Abh_reg[12] (.clk (\Clks[clk] ), .d (n_4239), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[12]));
  CDN_flop \Abh_reg[13] (.clk (\Clks[clk] ), .d (n_4240), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[13]));
  CDN_flop \Abh_reg[14] (.clk (\Clks[clk] ), .d (n_4241), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[14]));
  CDN_flop \Abh_reg[15] (.clk (\Clks[clk] ), .d (n_4242), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abh[15]));
  CDN_flop \Abl_reg[0] (.clk (\Clks[clk] ), .d (Abl[0]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[0]));
  CDN_flop \Abl_reg[1] (.clk (\Clks[clk] ), .d (Abl[1]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[1]));
  CDN_flop \Abl_reg[2] (.clk (\Clks[clk] ), .d (Abl[2]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[2]));
  CDN_flop \Abl_reg[3] (.clk (\Clks[clk] ), .d (Abl[3]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[3]));
  CDN_flop \Abl_reg[4] (.clk (\Clks[clk] ), .d (Abl[4]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[4]));
  CDN_flop \Abl_reg[5] (.clk (\Clks[clk] ), .d (Abl[5]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[5]));
  CDN_flop \Abl_reg[6] (.clk (\Clks[clk] ), .d (Abl[6]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[6]));
  CDN_flop \Abl_reg[7] (.clk (\Clks[clk] ), .d (Abl[7]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[7]));
  CDN_flop \Abl_reg[8] (.clk (\Clks[clk] ), .d (Abl[8]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[8]));
  CDN_flop \Abl_reg[9] (.clk (\Clks[clk] ), .d (Abl[9]), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[9]));
  CDN_flop \Abl_reg[10] (.clk (\Clks[clk] ), .d (Abl[10]), .sena
       (enT2), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[10]));
  CDN_flop \Abl_reg[11] (.clk (\Clks[clk] ), .d (Abl[11]), .sena
       (enT2), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[11]));
  CDN_flop \Abl_reg[12] (.clk (\Clks[clk] ), .d (Abl[12]), .sena
       (enT2), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[12]));
  CDN_flop \Abl_reg[13] (.clk (\Clks[clk] ), .d (Abl[13]), .sena
       (enT2), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[13]));
  CDN_flop \Abl_reg[14] (.clk (\Clks[clk] ), .d (Abl[14]), .sena
       (enT2), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[14]));
  CDN_flop \Abl_reg[15] (.clk (\Clks[clk] ), .d (Abl[15]), .sena
       (enT2), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (AblOut[15]));
  CDN_flop \Abd_reg[0] (.clk (\Clks[clk] ), .d (n_4243), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dcrInput[0]));
  CDN_flop \Abd_reg[1] (.clk (\Clks[clk] ), .d (n_4244), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dcrInput[1]));
  CDN_flop \Abd_reg[2] (.clk (\Clks[clk] ), .d (n_4245), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (dcrInput[2]));
  CDN_flop \Abd_reg[3] (.clk (\Clks[clk] ), .d (n_4246), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[3]));
  CDN_flop \Abd_reg[4] (.clk (\Clks[clk] ), .d (n_4247), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[4]));
  CDN_flop \Abd_reg[5] (.clk (\Clks[clk] ), .d (n_4248), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[5]));
  CDN_flop \Abd_reg[6] (.clk (\Clks[clk] ), .d (n_4249), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[6]));
  CDN_flop \Abd_reg[7] (.clk (\Clks[clk] ), .d (n_4250), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[7]));
  CDN_flop \Abd_reg[8] (.clk (\Clks[clk] ), .d (n_4251), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[8]));
  CDN_flop \Abd_reg[9] (.clk (\Clks[clk] ), .d (n_4252), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[9]));
  CDN_flop \Abd_reg[10] (.clk (\Clks[clk] ), .d (n_4253), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[10]));
  CDN_flop \Abd_reg[11] (.clk (\Clks[clk] ), .d (n_4254), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[11]));
  CDN_flop \Abd_reg[12] (.clk (\Clks[clk] ), .d (n_4255), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[12]));
  CDN_flop \Abd_reg[13] (.clk (\Clks[clk] ), .d (n_4256), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[13]));
  CDN_flop \Abd_reg[14] (.clk (\Clks[clk] ), .d (n_4257), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[14]));
  CDN_flop \Abd_reg[15] (.clk (\Clks[clk] ), .d (n_4258), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Abd[15]));
  CDN_flop \Dbd_reg[0] (.clk (\Clks[clk] ), .d (n_4259), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[0]));
  CDN_flop \Dbd_reg[1] (.clk (\Clks[clk] ), .d (n_4260), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[1]));
  CDN_flop \Dbd_reg[2] (.clk (\Clks[clk] ), .d (n_4261), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[2]));
  CDN_flop \Dbd_reg[3] (.clk (\Clks[clk] ), .d (n_4262), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[3]));
  CDN_flop \Dbd_reg[4] (.clk (\Clks[clk] ), .d (n_4263), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[4]));
  CDN_flop \Dbd_reg[5] (.clk (\Clks[clk] ), .d (n_4264), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[5]));
  CDN_flop \Dbd_reg[6] (.clk (\Clks[clk] ), .d (n_4265), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[6]));
  CDN_flop \Dbd_reg[7] (.clk (\Clks[clk] ), .d (n_4266), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[7]));
  CDN_flop \Dbd_reg[8] (.clk (\Clks[clk] ), .d (n_4267), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[8]));
  CDN_flop \Dbd_reg[9] (.clk (\Clks[clk] ), .d (n_4268), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[9]));
  CDN_flop \Dbd_reg[10] (.clk (\Clks[clk] ), .d (n_4269), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[10]));
  CDN_flop \Dbd_reg[11] (.clk (\Clks[clk] ), .d (n_4270), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[11]));
  CDN_flop \Dbd_reg[12] (.clk (\Clks[clk] ), .d (n_4271), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[12]));
  CDN_flop \Dbd_reg[13] (.clk (\Clks[clk] ), .d (n_4272), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[13]));
  CDN_flop \Dbd_reg[14] (.clk (\Clks[clk] ), .d (n_4273), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[14]));
  CDN_flop \Dbd_reg[15] (.clk (\Clks[clk] ), .d (n_4274), .sena (enT2),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (Dbd[15]));
  CDN_flop \preAbh_reg[0] (.clk (\Clks[clk] ), .d (abhMux[0]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[0]));
  CDN_flop \preAbh_reg[1] (.clk (\Clks[clk] ), .d (abhMux[1]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[1]));
  CDN_flop \preAbh_reg[2] (.clk (\Clks[clk] ), .d (abhMux[2]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[2]));
  CDN_flop \preAbh_reg[3] (.clk (\Clks[clk] ), .d (abhMux[3]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[3]));
  CDN_flop \preAbh_reg[4] (.clk (\Clks[clk] ), .d (abhMux[4]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[4]));
  CDN_flop \preAbh_reg[5] (.clk (\Clks[clk] ), .d (abhMux[5]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[5]));
  CDN_flop \preAbh_reg[6] (.clk (\Clks[clk] ), .d (abhMux[6]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[6]));
  CDN_flop \preAbh_reg[7] (.clk (\Clks[clk] ), .d (abhMux[7]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[7]));
  CDN_flop \preAbh_reg[8] (.clk (\Clks[clk] ), .d (abhMux[8]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[8]));
  CDN_flop \preAbh_reg[9] (.clk (\Clks[clk] ), .d (abhMux[9]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[9]));
  CDN_flop \preAbh_reg[10] (.clk (\Clks[clk] ), .d (abhMux[10]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[10]));
  CDN_flop \preAbh_reg[11] (.clk (\Clks[clk] ), .d (abhMux[11]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[11]));
  CDN_flop \preAbh_reg[12] (.clk (\Clks[clk] ), .d (abhMux[12]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[12]));
  CDN_flop \preAbh_reg[13] (.clk (\Clks[clk] ), .d (abhMux[13]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[13]));
  CDN_flop \preAbh_reg[14] (.clk (\Clks[clk] ), .d (abhMux[14]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[14]));
  CDN_flop \preAbh_reg[15] (.clk (\Clks[clk] ), .d (abhMux[15]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbh[15]));
  CDN_flop \preAbl_reg[0] (.clk (\Clks[clk] ), .d (ablMux[0]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[0]));
  CDN_flop \preAbl_reg[1] (.clk (\Clks[clk] ), .d (ablMux[1]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[1]));
  CDN_flop \preAbl_reg[2] (.clk (\Clks[clk] ), .d (ablMux[2]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[2]));
  CDN_flop \preAbl_reg[3] (.clk (\Clks[clk] ), .d (ablMux[3]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[3]));
  CDN_flop \preAbl_reg[4] (.clk (\Clks[clk] ), .d (ablMux[4]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[4]));
  CDN_flop \preAbl_reg[5] (.clk (\Clks[clk] ), .d (ablMux[5]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[5]));
  CDN_flop \preAbl_reg[6] (.clk (\Clks[clk] ), .d (ablMux[6]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[6]));
  CDN_flop \preAbl_reg[7] (.clk (\Clks[clk] ), .d (ablMux[7]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[7]));
  CDN_flop \preAbl_reg[8] (.clk (\Clks[clk] ), .d (ablMux[8]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[8]));
  CDN_flop \preAbl_reg[9] (.clk (\Clks[clk] ), .d (ablMux[9]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[9]));
  CDN_flop \preAbl_reg[10] (.clk (\Clks[clk] ), .d (ablMux[10]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[10]));
  CDN_flop \preAbl_reg[11] (.clk (\Clks[clk] ), .d (ablMux[11]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[11]));
  CDN_flop \preAbl_reg[12] (.clk (\Clks[clk] ), .d (ablMux[12]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[12]));
  CDN_flop \preAbl_reg[13] (.clk (\Clks[clk] ), .d (ablMux[13]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[13]));
  CDN_flop \preAbl_reg[14] (.clk (\Clks[clk] ), .d (ablMux[14]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[14]));
  CDN_flop \preAbl_reg[15] (.clk (\Clks[clk] ), .d (ablMux[15]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbl[15]));
  CDN_flop \preAbd_reg[0] (.clk (\Clks[clk] ), .d (abdMux[0]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[0]));
  CDN_flop \preAbd_reg[1] (.clk (\Clks[clk] ), .d (abdMux[1]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[1]));
  CDN_flop \preAbd_reg[2] (.clk (\Clks[clk] ), .d (abdMux[2]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[2]));
  CDN_flop \preAbd_reg[3] (.clk (\Clks[clk] ), .d (abdMux[3]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[3]));
  CDN_flop \preAbd_reg[4] (.clk (\Clks[clk] ), .d (abdMux[4]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[4]));
  CDN_flop \preAbd_reg[5] (.clk (\Clks[clk] ), .d (abdMux[5]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[5]));
  CDN_flop \preAbd_reg[6] (.clk (\Clks[clk] ), .d (abdMux[6]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[6]));
  CDN_flop \preAbd_reg[7] (.clk (\Clks[clk] ), .d (abdMux[7]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[7]));
  CDN_flop \preAbd_reg[8] (.clk (\Clks[clk] ), .d (abdMux[8]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[8]));
  CDN_flop \preAbd_reg[9] (.clk (\Clks[clk] ), .d (abdMux[9]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[9]));
  CDN_flop \preAbd_reg[10] (.clk (\Clks[clk] ), .d (abdMux[10]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[10]));
  CDN_flop \preAbd_reg[11] (.clk (\Clks[clk] ), .d (abdMux[11]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[11]));
  CDN_flop \preAbd_reg[12] (.clk (\Clks[clk] ), .d (abdMux[12]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[12]));
  CDN_flop \preAbd_reg[13] (.clk (\Clks[clk] ), .d (abdMux[13]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[13]));
  CDN_flop \preAbd_reg[14] (.clk (\Clks[clk] ), .d (abdMux[14]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[14]));
  CDN_flop \preAbd_reg[15] (.clk (\Clks[clk] ), .d (abdMux[15]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preAbd[15]));
  CDN_flop \preDbh_reg[0] (.clk (\Clks[clk] ), .d (dbhMux[0]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[0]));
  CDN_flop \preDbh_reg[1] (.clk (\Clks[clk] ), .d (dbhMux[1]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[1]));
  CDN_flop \preDbh_reg[2] (.clk (\Clks[clk] ), .d (dbhMux[2]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[2]));
  CDN_flop \preDbh_reg[3] (.clk (\Clks[clk] ), .d (dbhMux[3]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[3]));
  CDN_flop \preDbh_reg[4] (.clk (\Clks[clk] ), .d (dbhMux[4]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[4]));
  CDN_flop \preDbh_reg[5] (.clk (\Clks[clk] ), .d (dbhMux[5]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[5]));
  CDN_flop \preDbh_reg[6] (.clk (\Clks[clk] ), .d (dbhMux[6]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[6]));
  CDN_flop \preDbh_reg[7] (.clk (\Clks[clk] ), .d (dbhMux[7]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[7]));
  CDN_flop \preDbh_reg[8] (.clk (\Clks[clk] ), .d (dbhMux[8]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[8]));
  CDN_flop \preDbh_reg[9] (.clk (\Clks[clk] ), .d (dbhMux[9]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[9]));
  CDN_flop \preDbh_reg[10] (.clk (\Clks[clk] ), .d (dbhMux[10]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[10]));
  CDN_flop \preDbh_reg[11] (.clk (\Clks[clk] ), .d (dbhMux[11]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[11]));
  CDN_flop \preDbh_reg[12] (.clk (\Clks[clk] ), .d (dbhMux[12]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[12]));
  CDN_flop \preDbh_reg[13] (.clk (\Clks[clk] ), .d (dbhMux[13]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[13]));
  CDN_flop \preDbh_reg[14] (.clk (\Clks[clk] ), .d (dbhMux[14]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[14]));
  CDN_flop \preDbh_reg[15] (.clk (\Clks[clk] ), .d (dbhMux[15]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbh[15]));
  CDN_flop \preDbl_reg[0] (.clk (\Clks[clk] ), .d (dblMux[0]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[0]));
  CDN_flop \preDbl_reg[1] (.clk (\Clks[clk] ), .d (dblMux[1]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[1]));
  CDN_flop \preDbl_reg[2] (.clk (\Clks[clk] ), .d (dblMux[2]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[2]));
  CDN_flop \preDbl_reg[3] (.clk (\Clks[clk] ), .d (dblMux[3]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[3]));
  CDN_flop \preDbl_reg[4] (.clk (\Clks[clk] ), .d (dblMux[4]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[4]));
  CDN_flop \preDbl_reg[5] (.clk (\Clks[clk] ), .d (dblMux[5]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[5]));
  CDN_flop \preDbl_reg[6] (.clk (\Clks[clk] ), .d (dblMux[6]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[6]));
  CDN_flop \preDbl_reg[7] (.clk (\Clks[clk] ), .d (dblMux[7]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[7]));
  CDN_flop \preDbl_reg[8] (.clk (\Clks[clk] ), .d (dblMux[8]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[8]));
  CDN_flop \preDbl_reg[9] (.clk (\Clks[clk] ), .d (dblMux[9]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[9]));
  CDN_flop \preDbl_reg[10] (.clk (\Clks[clk] ), .d (dblMux[10]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[10]));
  CDN_flop \preDbl_reg[11] (.clk (\Clks[clk] ), .d (dblMux[11]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[11]));
  CDN_flop \preDbl_reg[12] (.clk (\Clks[clk] ), .d (dblMux[12]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[12]));
  CDN_flop \preDbl_reg[13] (.clk (\Clks[clk] ), .d (dblMux[13]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[13]));
  CDN_flop \preDbl_reg[14] (.clk (\Clks[clk] ), .d (dblMux[14]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[14]));
  CDN_flop \preDbl_reg[15] (.clk (\Clks[clk] ), .d (dblMux[15]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbl[15]));
  CDN_flop \preDbd_reg[0] (.clk (\Clks[clk] ), .d (dbdMux[0]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[0]));
  CDN_flop \preDbd_reg[1] (.clk (\Clks[clk] ), .d (dbdMux[1]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[1]));
  CDN_flop \preDbd_reg[2] (.clk (\Clks[clk] ), .d (dbdMux[2]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[2]));
  CDN_flop \preDbd_reg[3] (.clk (\Clks[clk] ), .d (dbdMux[3]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[3]));
  CDN_flop \preDbd_reg[4] (.clk (\Clks[clk] ), .d (dbdMux[4]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[4]));
  CDN_flop \preDbd_reg[5] (.clk (\Clks[clk] ), .d (dbdMux[5]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[5]));
  CDN_flop \preDbd_reg[6] (.clk (\Clks[clk] ), .d (dbdMux[6]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[6]));
  CDN_flop \preDbd_reg[7] (.clk (\Clks[clk] ), .d (dbdMux[7]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[7]));
  CDN_flop \preDbd_reg[8] (.clk (\Clks[clk] ), .d (dbdMux[8]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[8]));
  CDN_flop \preDbd_reg[9] (.clk (\Clks[clk] ), .d (dbdMux[9]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[9]));
  CDN_flop \preDbd_reg[10] (.clk (\Clks[clk] ), .d (dbdMux[10]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[10]));
  CDN_flop \preDbd_reg[11] (.clk (\Clks[clk] ), .d (dbdMux[11]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[11]));
  CDN_flop \preDbd_reg[12] (.clk (\Clks[clk] ), .d (dbdMux[12]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[12]));
  CDN_flop \preDbd_reg[13] (.clk (\Clks[clk] ), .d (dbdMux[13]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[13]));
  CDN_flop \preDbd_reg[14] (.clk (\Clks[clk] ), .d (dbdMux[14]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[14]));
  CDN_flop \preDbd_reg[15] (.clk (\Clks[clk] ), .d (dbdMux[15]), .sena
       (enT1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (preDbd[15]));
  CDN_flop \aob_reg[0] (.clk (\Clks[clk] ), .d (n_4282), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob0));
  CDN_flop \aob_reg[1] (.clk (\Clks[clk] ), .d (n_4284), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[1]));
  CDN_flop \aob_reg[2] (.clk (\Clks[clk] ), .d (n_4285), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[2]));
  CDN_flop \aob_reg[3] (.clk (\Clks[clk] ), .d (n_4286), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[3]));
  CDN_flop \aob_reg[4] (.clk (\Clks[clk] ), .d (n_4287), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[4]));
  CDN_flop \aob_reg[5] (.clk (\Clks[clk] ), .d (n_4288), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[5]));
  CDN_flop \aob_reg[6] (.clk (\Clks[clk] ), .d (n_4289), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[6]));
  CDN_flop \aob_reg[7] (.clk (\Clks[clk] ), .d (n_4290), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[7]));
  CDN_flop \aob_reg[8] (.clk (\Clks[clk] ), .d (n_4291), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[8]));
  CDN_flop \aob_reg[9] (.clk (\Clks[clk] ), .d (n_4292), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[9]));
  CDN_flop \aob_reg[10] (.clk (\Clks[clk] ), .d (n_4293), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[10]));
  CDN_flop \aob_reg[11] (.clk (\Clks[clk] ), .d (n_4294), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[11]));
  CDN_flop \aob_reg[12] (.clk (\Clks[clk] ), .d (n_4295), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[12]));
  CDN_flop \aob_reg[13] (.clk (\Clks[clk] ), .d (n_4296), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[13]));
  CDN_flop \aob_reg[14] (.clk (\Clks[clk] ), .d (n_4297), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[14]));
  CDN_flop \aob_reg[15] (.clk (\Clks[clk] ), .d (n_4298), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[15]));
  CDN_flop \aob_reg[16] (.clk (\Clks[clk] ), .d (n_4299), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[16]));
  CDN_flop \aob_reg[17] (.clk (\Clks[clk] ), .d (n_4300), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[17]));
  CDN_flop \aob_reg[18] (.clk (\Clks[clk] ), .d (n_4301), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[18]));
  CDN_flop \aob_reg[19] (.clk (\Clks[clk] ), .d (n_4302), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[19]));
  CDN_flop \aob_reg[20] (.clk (\Clks[clk] ), .d (n_4303), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[20]));
  CDN_flop \aob_reg[21] (.clk (\Clks[clk] ), .d (n_4304), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[21]));
  CDN_flop \aob_reg[22] (.clk (\Clks[clk] ), .d (n_4305), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[22]));
  CDN_flop \aob_reg[23] (.clk (\Clks[clk] ), .d (n_4306), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (eab[23]));
  CDN_flop \aob_reg[24] (.clk (\Clks[clk] ), .d (n_4307), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[24]));
  CDN_flop \aob_reg[25] (.clk (\Clks[clk] ), .d (n_4308), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[25]));
  CDN_flop \aob_reg[26] (.clk (\Clks[clk] ), .d (n_4309), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[26]));
  CDN_flop \aob_reg[27] (.clk (\Clks[clk] ), .d (n_4310), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[27]));
  CDN_flop \aob_reg[28] (.clk (\Clks[clk] ), .d (n_4311), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[28]));
  CDN_flop \aob_reg[29] (.clk (\Clks[clk] ), .d (n_4312), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[29]));
  CDN_flop \aob_reg[30] (.clk (\Clks[clk] ), .d (n_4313), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[30]));
  CDN_flop \aob_reg[31] (.clk (\Clks[clk] ), .d (n_4314), .sena
       (n_4283), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (aob[31]));
  CDN_flop \auReg_reg[0] (.clk (\Clks[clk] ), .d (n_1234), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[0]));
  CDN_flop \auReg_reg[1] (.clk (\Clks[clk] ), .d (n_1235), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[1]));
  CDN_flop \auReg_reg[2] (.clk (\Clks[clk] ), .d (n_1236), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[2]));
  CDN_flop \auReg_reg[3] (.clk (\Clks[clk] ), .d (n_1237), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[3]));
  CDN_flop \auReg_reg[4] (.clk (\Clks[clk] ), .d (n_1238), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[4]));
  CDN_flop \auReg_reg[5] (.clk (\Clks[clk] ), .d (n_1239), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[5]));
  CDN_flop \auReg_reg[6] (.clk (\Clks[clk] ), .d (n_1240), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[6]));
  CDN_flop \auReg_reg[7] (.clk (\Clks[clk] ), .d (n_1241), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[7]));
  CDN_flop \auReg_reg[8] (.clk (\Clks[clk] ), .d (n_1242), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[8]));
  CDN_flop \auReg_reg[9] (.clk (\Clks[clk] ), .d (n_1243), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[9]));
  CDN_flop \auReg_reg[10] (.clk (\Clks[clk] ), .d (n_1244), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[10]));
  CDN_flop \auReg_reg[11] (.clk (\Clks[clk] ), .d (n_1245), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[11]));
  CDN_flop \auReg_reg[12] (.clk (\Clks[clk] ), .d (n_1246), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[12]));
  CDN_flop \auReg_reg[13] (.clk (\Clks[clk] ), .d (n_1247), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[13]));
  CDN_flop \auReg_reg[14] (.clk (\Clks[clk] ), .d (n_1248), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[14]));
  CDN_flop \auReg_reg[15] (.clk (\Clks[clk] ), .d (n_1249), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[15]));
  CDN_flop \auReg_reg[16] (.clk (\Clks[clk] ), .d (n_1250), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[16]));
  CDN_flop \auReg_reg[17] (.clk (\Clks[clk] ), .d (n_1251), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[17]));
  CDN_flop \auReg_reg[18] (.clk (\Clks[clk] ), .d (n_1252), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[18]));
  CDN_flop \auReg_reg[19] (.clk (\Clks[clk] ), .d (n_1253), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[19]));
  CDN_flop \auReg_reg[20] (.clk (\Clks[clk] ), .d (n_1254), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[20]));
  CDN_flop \auReg_reg[21] (.clk (\Clks[clk] ), .d (n_1255), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[21]));
  CDN_flop \auReg_reg[22] (.clk (\Clks[clk] ), .d (n_1256), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[22]));
  CDN_flop \auReg_reg[23] (.clk (\Clks[clk] ), .d (n_1257), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[23]));
  CDN_flop \auReg_reg[24] (.clk (\Clks[clk] ), .d (n_1258), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[24]));
  CDN_flop \auReg_reg[25] (.clk (\Clks[clk] ), .d (n_1259), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[25]));
  CDN_flop \auReg_reg[26] (.clk (\Clks[clk] ), .d (n_1260), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[26]));
  CDN_flop \auReg_reg[27] (.clk (\Clks[clk] ), .d (n_1261), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[27]));
  CDN_flop \auReg_reg[28] (.clk (\Clks[clk] ), .d (n_1262), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[28]));
  CDN_flop \auReg_reg[29] (.clk (\Clks[clk] ), .d (n_1263), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[29]));
  CDN_flop \auReg_reg[30] (.clk (\Clks[clk] ), .d (n_1264), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[30]));
  CDN_flop \auReg_reg[31] (.clk (\Clks[clk] ), .d (n_1265), .sena
       (n_453), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (auReg[31]));
  CDN_flop \regs68L_reg[17][0] (.clk (\Clks[clk] ), .d (n_4382), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [0]));
  CDN_flop \regs68L_reg[17][1] (.clk (\Clks[clk] ), .d (n_4384), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [1]));
  CDN_flop \regs68L_reg[17][2] (.clk (\Clks[clk] ), .d (n_4385), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [2]));
  CDN_flop \regs68L_reg[17][3] (.clk (\Clks[clk] ), .d (n_4386), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [3]));
  CDN_flop \regs68L_reg[17][4] (.clk (\Clks[clk] ), .d (n_4387), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [4]));
  CDN_flop \regs68L_reg[17][5] (.clk (\Clks[clk] ), .d (n_4388), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [5]));
  CDN_flop \regs68L_reg[17][6] (.clk (\Clks[clk] ), .d (n_4389), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [6]));
  CDN_flop \regs68L_reg[17][7] (.clk (\Clks[clk] ), .d (n_4390), .sena
       (n_4383), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [7]));
  CDN_flop \regs68L_reg[17][8] (.clk (\Clks[clk] ), .d (n_4391), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [8]));
  CDN_flop \regs68L_reg[17][9] (.clk (\Clks[clk] ), .d (n_4393), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [9]));
  CDN_flop \regs68L_reg[17][10] (.clk (\Clks[clk] ), .d (n_4394), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [10]));
  CDN_flop \regs68L_reg[17][11] (.clk (\Clks[clk] ), .d (n_4395), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [11]));
  CDN_flop \regs68L_reg[17][12] (.clk (\Clks[clk] ), .d (n_4396), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [12]));
  CDN_flop \regs68L_reg[17][13] (.clk (\Clks[clk] ), .d (n_4397), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [13]));
  CDN_flop \regs68L_reg[17][14] (.clk (\Clks[clk] ), .d (n_4398), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [14]));
  CDN_flop \regs68L_reg[17][15] (.clk (\Clks[clk] ), .d (n_4399), .sena
       (n_4392), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[17] [15]));
  CDN_flop \regs68L_reg[16][0] (.clk (\Clks[clk] ), .d (n_4461), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [0]));
  CDN_flop \regs68L_reg[16][1] (.clk (\Clks[clk] ), .d (n_4463), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [1]));
  CDN_flop \regs68L_reg[16][2] (.clk (\Clks[clk] ), .d (n_4464), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [2]));
  CDN_flop \regs68L_reg[16][3] (.clk (\Clks[clk] ), .d (n_4465), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [3]));
  CDN_flop \regs68L_reg[16][4] (.clk (\Clks[clk] ), .d (n_4466), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [4]));
  CDN_flop \regs68L_reg[16][5] (.clk (\Clks[clk] ), .d (n_4467), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [5]));
  CDN_flop \regs68L_reg[16][6] (.clk (\Clks[clk] ), .d (n_4468), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [6]));
  CDN_flop \regs68L_reg[16][7] (.clk (\Clks[clk] ), .d (n_4469), .sena
       (n_4462), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [7]));
  CDN_flop \regs68L_reg[16][8] (.clk (\Clks[clk] ), .d (n_4470), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [8]));
  CDN_flop \regs68L_reg[16][9] (.clk (\Clks[clk] ), .d (n_4472), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [9]));
  CDN_flop \regs68L_reg[16][10] (.clk (\Clks[clk] ), .d (n_4473), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [10]));
  CDN_flop \regs68L_reg[16][11] (.clk (\Clks[clk] ), .d (n_4474), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [11]));
  CDN_flop \regs68L_reg[16][12] (.clk (\Clks[clk] ), .d (n_4475), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [12]));
  CDN_flop \regs68L_reg[16][13] (.clk (\Clks[clk] ), .d (n_4476), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [13]));
  CDN_flop \regs68L_reg[16][14] (.clk (\Clks[clk] ), .d (n_4477), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [14]));
  CDN_flop \regs68L_reg[16][15] (.clk (\Clks[clk] ), .d (n_4478), .sena
       (n_4471), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[16] [15]));
  CDN_flop \regs68L_reg[15][0] (.clk (\Clks[clk] ), .d (n_4540), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [0]));
  CDN_flop \regs68L_reg[15][1] (.clk (\Clks[clk] ), .d (n_4542), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [1]));
  CDN_flop \regs68L_reg[15][2] (.clk (\Clks[clk] ), .d (n_4543), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [2]));
  CDN_flop \regs68L_reg[15][3] (.clk (\Clks[clk] ), .d (n_4544), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [3]));
  CDN_flop \regs68L_reg[15][4] (.clk (\Clks[clk] ), .d (n_4545), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [4]));
  CDN_flop \regs68L_reg[15][5] (.clk (\Clks[clk] ), .d (n_4546), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [5]));
  CDN_flop \regs68L_reg[15][6] (.clk (\Clks[clk] ), .d (n_4547), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [6]));
  CDN_flop \regs68L_reg[15][7] (.clk (\Clks[clk] ), .d (n_4548), .sena
       (n_4541), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [7]));
  CDN_flop \regs68L_reg[15][8] (.clk (\Clks[clk] ), .d (n_4549), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [8]));
  CDN_flop \regs68L_reg[15][9] (.clk (\Clks[clk] ), .d (n_4551), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [9]));
  CDN_flop \regs68L_reg[15][10] (.clk (\Clks[clk] ), .d (n_4552), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [10]));
  CDN_flop \regs68L_reg[15][11] (.clk (\Clks[clk] ), .d (n_4553), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [11]));
  CDN_flop \regs68L_reg[15][12] (.clk (\Clks[clk] ), .d (n_4554), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [12]));
  CDN_flop \regs68L_reg[15][13] (.clk (\Clks[clk] ), .d (n_4555), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [13]));
  CDN_flop \regs68L_reg[15][14] (.clk (\Clks[clk] ), .d (n_4556), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [14]));
  CDN_flop \regs68L_reg[15][15] (.clk (\Clks[clk] ), .d (n_4557), .sena
       (n_4550), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[15] [15]));
  CDN_flop \regs68L_reg[14][0] (.clk (\Clks[clk] ), .d (n_4619), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [0]));
  CDN_flop \regs68L_reg[14][1] (.clk (\Clks[clk] ), .d (n_4621), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [1]));
  CDN_flop \regs68L_reg[14][2] (.clk (\Clks[clk] ), .d (n_4622), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [2]));
  CDN_flop \regs68L_reg[14][3] (.clk (\Clks[clk] ), .d (n_4623), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [3]));
  CDN_flop \regs68L_reg[14][4] (.clk (\Clks[clk] ), .d (n_4624), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [4]));
  CDN_flop \regs68L_reg[14][5] (.clk (\Clks[clk] ), .d (n_4625), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [5]));
  CDN_flop \regs68L_reg[14][6] (.clk (\Clks[clk] ), .d (n_4626), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [6]));
  CDN_flop \regs68L_reg[14][7] (.clk (\Clks[clk] ), .d (n_4627), .sena
       (n_4620), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [7]));
  CDN_flop \regs68L_reg[14][8] (.clk (\Clks[clk] ), .d (n_4628), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [8]));
  CDN_flop \regs68L_reg[14][9] (.clk (\Clks[clk] ), .d (n_4630), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [9]));
  CDN_flop \regs68L_reg[14][10] (.clk (\Clks[clk] ), .d (n_4631), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [10]));
  CDN_flop \regs68L_reg[14][11] (.clk (\Clks[clk] ), .d (n_4632), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [11]));
  CDN_flop \regs68L_reg[14][12] (.clk (\Clks[clk] ), .d (n_4633), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [12]));
  CDN_flop \regs68L_reg[14][13] (.clk (\Clks[clk] ), .d (n_4634), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [13]));
  CDN_flop \regs68L_reg[14][14] (.clk (\Clks[clk] ), .d (n_4635), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [14]));
  CDN_flop \regs68L_reg[14][15] (.clk (\Clks[clk] ), .d (n_4636), .sena
       (n_4629), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[14] [15]));
  CDN_flop \regs68L_reg[13][0] (.clk (\Clks[clk] ), .d (n_4698), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [0]));
  CDN_flop \regs68L_reg[13][1] (.clk (\Clks[clk] ), .d (n_4700), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [1]));
  CDN_flop \regs68L_reg[13][2] (.clk (\Clks[clk] ), .d (n_4701), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [2]));
  CDN_flop \regs68L_reg[13][3] (.clk (\Clks[clk] ), .d (n_4702), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [3]));
  CDN_flop \regs68L_reg[13][4] (.clk (\Clks[clk] ), .d (n_4703), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [4]));
  CDN_flop \regs68L_reg[13][5] (.clk (\Clks[clk] ), .d (n_4704), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [5]));
  CDN_flop \regs68L_reg[13][6] (.clk (\Clks[clk] ), .d (n_4705), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [6]));
  CDN_flop \regs68L_reg[13][7] (.clk (\Clks[clk] ), .d (n_4706), .sena
       (n_4699), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [7]));
  CDN_flop \regs68L_reg[13][8] (.clk (\Clks[clk] ), .d (n_4707), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [8]));
  CDN_flop \regs68L_reg[13][9] (.clk (\Clks[clk] ), .d (n_4709), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [9]));
  CDN_flop \regs68L_reg[13][10] (.clk (\Clks[clk] ), .d (n_4710), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [10]));
  CDN_flop \regs68L_reg[13][11] (.clk (\Clks[clk] ), .d (n_4711), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [11]));
  CDN_flop \regs68L_reg[13][12] (.clk (\Clks[clk] ), .d (n_4712), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [12]));
  CDN_flop \regs68L_reg[13][13] (.clk (\Clks[clk] ), .d (n_4713), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [13]));
  CDN_flop \regs68L_reg[13][14] (.clk (\Clks[clk] ), .d (n_4714), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [14]));
  CDN_flop \regs68L_reg[13][15] (.clk (\Clks[clk] ), .d (n_4715), .sena
       (n_4708), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[13] [15]));
  CDN_flop \regs68L_reg[12][0] (.clk (\Clks[clk] ), .d (n_4777), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [0]));
  CDN_flop \regs68L_reg[12][1] (.clk (\Clks[clk] ), .d (n_4779), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [1]));
  CDN_flop \regs68L_reg[12][2] (.clk (\Clks[clk] ), .d (n_4780), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [2]));
  CDN_flop \regs68L_reg[12][3] (.clk (\Clks[clk] ), .d (n_4781), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [3]));
  CDN_flop \regs68L_reg[12][4] (.clk (\Clks[clk] ), .d (n_4782), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [4]));
  CDN_flop \regs68L_reg[12][5] (.clk (\Clks[clk] ), .d (n_4783), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [5]));
  CDN_flop \regs68L_reg[12][6] (.clk (\Clks[clk] ), .d (n_4784), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [6]));
  CDN_flop \regs68L_reg[12][7] (.clk (\Clks[clk] ), .d (n_4785), .sena
       (n_4778), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [7]));
  CDN_flop \regs68L_reg[12][8] (.clk (\Clks[clk] ), .d (n_4786), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [8]));
  CDN_flop \regs68L_reg[12][9] (.clk (\Clks[clk] ), .d (n_4788), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [9]));
  CDN_flop \regs68L_reg[12][10] (.clk (\Clks[clk] ), .d (n_4789), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [10]));
  CDN_flop \regs68L_reg[12][11] (.clk (\Clks[clk] ), .d (n_4790), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [11]));
  CDN_flop \regs68L_reg[12][12] (.clk (\Clks[clk] ), .d (n_4791), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [12]));
  CDN_flop \regs68L_reg[12][13] (.clk (\Clks[clk] ), .d (n_4792), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [13]));
  CDN_flop \regs68L_reg[12][14] (.clk (\Clks[clk] ), .d (n_4793), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [14]));
  CDN_flop \regs68L_reg[12][15] (.clk (\Clks[clk] ), .d (n_4794), .sena
       (n_4787), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[12] [15]));
  CDN_flop \regs68L_reg[11][0] (.clk (\Clks[clk] ), .d (n_4856), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [0]));
  CDN_flop \regs68L_reg[11][1] (.clk (\Clks[clk] ), .d (n_4858), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [1]));
  CDN_flop \regs68L_reg[11][2] (.clk (\Clks[clk] ), .d (n_4859), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [2]));
  CDN_flop \regs68L_reg[11][3] (.clk (\Clks[clk] ), .d (n_4860), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [3]));
  CDN_flop \regs68L_reg[11][4] (.clk (\Clks[clk] ), .d (n_4861), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [4]));
  CDN_flop \regs68L_reg[11][5] (.clk (\Clks[clk] ), .d (n_4862), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [5]));
  CDN_flop \regs68L_reg[11][6] (.clk (\Clks[clk] ), .d (n_4863), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [6]));
  CDN_flop \regs68L_reg[11][7] (.clk (\Clks[clk] ), .d (n_4864), .sena
       (n_4857), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [7]));
  CDN_flop \regs68L_reg[11][8] (.clk (\Clks[clk] ), .d (n_4865), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [8]));
  CDN_flop \regs68L_reg[11][9] (.clk (\Clks[clk] ), .d (n_4867), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [9]));
  CDN_flop \regs68L_reg[11][10] (.clk (\Clks[clk] ), .d (n_4868), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [10]));
  CDN_flop \regs68L_reg[11][11] (.clk (\Clks[clk] ), .d (n_4869), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [11]));
  CDN_flop \regs68L_reg[11][12] (.clk (\Clks[clk] ), .d (n_4870), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [12]));
  CDN_flop \regs68L_reg[11][13] (.clk (\Clks[clk] ), .d (n_4871), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [13]));
  CDN_flop \regs68L_reg[11][14] (.clk (\Clks[clk] ), .d (n_4872), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [14]));
  CDN_flop \regs68L_reg[11][15] (.clk (\Clks[clk] ), .d (n_4873), .sena
       (n_4866), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[11] [15]));
  CDN_flop \regs68L_reg[10][0] (.clk (\Clks[clk] ), .d (n_4935), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [0]));
  CDN_flop \regs68L_reg[10][1] (.clk (\Clks[clk] ), .d (n_4937), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [1]));
  CDN_flop \regs68L_reg[10][2] (.clk (\Clks[clk] ), .d (n_4938), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [2]));
  CDN_flop \regs68L_reg[10][3] (.clk (\Clks[clk] ), .d (n_4939), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [3]));
  CDN_flop \regs68L_reg[10][4] (.clk (\Clks[clk] ), .d (n_4940), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [4]));
  CDN_flop \regs68L_reg[10][5] (.clk (\Clks[clk] ), .d (n_4941), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [5]));
  CDN_flop \regs68L_reg[10][6] (.clk (\Clks[clk] ), .d (n_4942), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [6]));
  CDN_flop \regs68L_reg[10][7] (.clk (\Clks[clk] ), .d (n_4943), .sena
       (n_4936), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [7]));
  CDN_flop \regs68L_reg[10][8] (.clk (\Clks[clk] ), .d (n_4944), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [8]));
  CDN_flop \regs68L_reg[10][9] (.clk (\Clks[clk] ), .d (n_4946), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [9]));
  CDN_flop \regs68L_reg[10][10] (.clk (\Clks[clk] ), .d (n_4947), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [10]));
  CDN_flop \regs68L_reg[10][11] (.clk (\Clks[clk] ), .d (n_4948), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [11]));
  CDN_flop \regs68L_reg[10][12] (.clk (\Clks[clk] ), .d (n_4949), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [12]));
  CDN_flop \regs68L_reg[10][13] (.clk (\Clks[clk] ), .d (n_4950), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [13]));
  CDN_flop \regs68L_reg[10][14] (.clk (\Clks[clk] ), .d (n_4951), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [14]));
  CDN_flop \regs68L_reg[10][15] (.clk (\Clks[clk] ), .d (n_4952), .sena
       (n_4945), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[10] [15]));
  CDN_flop \regs68L_reg[9][0] (.clk (\Clks[clk] ), .d (n_5014), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [0]));
  CDN_flop \regs68L_reg[9][1] (.clk (\Clks[clk] ), .d (n_5016), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [1]));
  CDN_flop \regs68L_reg[9][2] (.clk (\Clks[clk] ), .d (n_5017), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [2]));
  CDN_flop \regs68L_reg[9][3] (.clk (\Clks[clk] ), .d (n_5018), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [3]));
  CDN_flop \regs68L_reg[9][4] (.clk (\Clks[clk] ), .d (n_5019), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [4]));
  CDN_flop \regs68L_reg[9][5] (.clk (\Clks[clk] ), .d (n_5020), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [5]));
  CDN_flop \regs68L_reg[9][6] (.clk (\Clks[clk] ), .d (n_5021), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [6]));
  CDN_flop \regs68L_reg[9][7] (.clk (\Clks[clk] ), .d (n_5022), .sena
       (n_5015), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [7]));
  CDN_flop \regs68L_reg[9][8] (.clk (\Clks[clk] ), .d (n_5023), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [8]));
  CDN_flop \regs68L_reg[9][9] (.clk (\Clks[clk] ), .d (n_5025), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [9]));
  CDN_flop \regs68L_reg[9][10] (.clk (\Clks[clk] ), .d (n_5026), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [10]));
  CDN_flop \regs68L_reg[9][11] (.clk (\Clks[clk] ), .d (n_5027), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [11]));
  CDN_flop \regs68L_reg[9][12] (.clk (\Clks[clk] ), .d (n_5028), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [12]));
  CDN_flop \regs68L_reg[9][13] (.clk (\Clks[clk] ), .d (n_5029), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [13]));
  CDN_flop \regs68L_reg[9][14] (.clk (\Clks[clk] ), .d (n_5030), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [14]));
  CDN_flop \regs68L_reg[9][15] (.clk (\Clks[clk] ), .d (n_5031), .sena
       (n_5024), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[9] [15]));
  CDN_flop \regs68L_reg[8][0] (.clk (\Clks[clk] ), .d (n_5093), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [0]));
  CDN_flop \regs68L_reg[8][1] (.clk (\Clks[clk] ), .d (n_5095), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [1]));
  CDN_flop \regs68L_reg[8][2] (.clk (\Clks[clk] ), .d (n_5096), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [2]));
  CDN_flop \regs68L_reg[8][3] (.clk (\Clks[clk] ), .d (n_5097), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [3]));
  CDN_flop \regs68L_reg[8][4] (.clk (\Clks[clk] ), .d (n_5098), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [4]));
  CDN_flop \regs68L_reg[8][5] (.clk (\Clks[clk] ), .d (n_5099), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [5]));
  CDN_flop \regs68L_reg[8][6] (.clk (\Clks[clk] ), .d (n_5100), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [6]));
  CDN_flop \regs68L_reg[8][7] (.clk (\Clks[clk] ), .d (n_5101), .sena
       (n_5094), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [7]));
  CDN_flop \regs68L_reg[8][8] (.clk (\Clks[clk] ), .d (n_5102), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [8]));
  CDN_flop \regs68L_reg[8][9] (.clk (\Clks[clk] ), .d (n_5104), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [9]));
  CDN_flop \regs68L_reg[8][10] (.clk (\Clks[clk] ), .d (n_5105), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [10]));
  CDN_flop \regs68L_reg[8][11] (.clk (\Clks[clk] ), .d (n_5106), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [11]));
  CDN_flop \regs68L_reg[8][12] (.clk (\Clks[clk] ), .d (n_5107), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [12]));
  CDN_flop \regs68L_reg[8][13] (.clk (\Clks[clk] ), .d (n_5108), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [13]));
  CDN_flop \regs68L_reg[8][14] (.clk (\Clks[clk] ), .d (n_5109), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [14]));
  CDN_flop \regs68L_reg[8][15] (.clk (\Clks[clk] ), .d (n_5110), .sena
       (n_5103), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[8] [15]));
  CDN_flop \regs68L_reg[7][0] (.clk (\Clks[clk] ), .d (n_5172), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [0]));
  CDN_flop \regs68L_reg[7][1] (.clk (\Clks[clk] ), .d (n_5174), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [1]));
  CDN_flop \regs68L_reg[7][2] (.clk (\Clks[clk] ), .d (n_5175), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [2]));
  CDN_flop \regs68L_reg[7][3] (.clk (\Clks[clk] ), .d (n_5176), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [3]));
  CDN_flop \regs68L_reg[7][4] (.clk (\Clks[clk] ), .d (n_5177), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [4]));
  CDN_flop \regs68L_reg[7][5] (.clk (\Clks[clk] ), .d (n_5178), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [5]));
  CDN_flop \regs68L_reg[7][6] (.clk (\Clks[clk] ), .d (n_5179), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [6]));
  CDN_flop \regs68L_reg[7][7] (.clk (\Clks[clk] ), .d (n_5180), .sena
       (n_5173), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [7]));
  CDN_flop \regs68L_reg[7][8] (.clk (\Clks[clk] ), .d (n_5181), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [8]));
  CDN_flop \regs68L_reg[7][9] (.clk (\Clks[clk] ), .d (n_5183), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [9]));
  CDN_flop \regs68L_reg[7][10] (.clk (\Clks[clk] ), .d (n_5184), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [10]));
  CDN_flop \regs68L_reg[7][11] (.clk (\Clks[clk] ), .d (n_5185), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [11]));
  CDN_flop \regs68L_reg[7][12] (.clk (\Clks[clk] ), .d (n_5186), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [12]));
  CDN_flop \regs68L_reg[7][13] (.clk (\Clks[clk] ), .d (n_5187), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [13]));
  CDN_flop \regs68L_reg[7][14] (.clk (\Clks[clk] ), .d (n_5188), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [14]));
  CDN_flop \regs68L_reg[7][15] (.clk (\Clks[clk] ), .d (n_5189), .sena
       (n_5182), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[7] [15]));
  CDN_flop \regs68L_reg[6][0] (.clk (\Clks[clk] ), .d (n_5251), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [0]));
  CDN_flop \regs68L_reg[6][1] (.clk (\Clks[clk] ), .d (n_5253), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [1]));
  CDN_flop \regs68L_reg[6][2] (.clk (\Clks[clk] ), .d (n_5254), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [2]));
  CDN_flop \regs68L_reg[6][3] (.clk (\Clks[clk] ), .d (n_5255), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [3]));
  CDN_flop \regs68L_reg[6][4] (.clk (\Clks[clk] ), .d (n_5256), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [4]));
  CDN_flop \regs68L_reg[6][5] (.clk (\Clks[clk] ), .d (n_5257), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [5]));
  CDN_flop \regs68L_reg[6][6] (.clk (\Clks[clk] ), .d (n_5258), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [6]));
  CDN_flop \regs68L_reg[6][7] (.clk (\Clks[clk] ), .d (n_5259), .sena
       (n_5252), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [7]));
  CDN_flop \regs68L_reg[6][8] (.clk (\Clks[clk] ), .d (n_5260), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [8]));
  CDN_flop \regs68L_reg[6][9] (.clk (\Clks[clk] ), .d (n_5262), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [9]));
  CDN_flop \regs68L_reg[6][10] (.clk (\Clks[clk] ), .d (n_5263), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [10]));
  CDN_flop \regs68L_reg[6][11] (.clk (\Clks[clk] ), .d (n_5264), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [11]));
  CDN_flop \regs68L_reg[6][12] (.clk (\Clks[clk] ), .d (n_5265), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [12]));
  CDN_flop \regs68L_reg[6][13] (.clk (\Clks[clk] ), .d (n_5266), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [13]));
  CDN_flop \regs68L_reg[6][14] (.clk (\Clks[clk] ), .d (n_5267), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [14]));
  CDN_flop \regs68L_reg[6][15] (.clk (\Clks[clk] ), .d (n_5268), .sena
       (n_5261), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[6] [15]));
  CDN_flop \regs68L_reg[5][0] (.clk (\Clks[clk] ), .d (n_5330), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [0]));
  CDN_flop \regs68L_reg[5][1] (.clk (\Clks[clk] ), .d (n_5332), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [1]));
  CDN_flop \regs68L_reg[5][2] (.clk (\Clks[clk] ), .d (n_5333), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [2]));
  CDN_flop \regs68L_reg[5][3] (.clk (\Clks[clk] ), .d (n_5334), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [3]));
  CDN_flop \regs68L_reg[5][4] (.clk (\Clks[clk] ), .d (n_5335), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [4]));
  CDN_flop \regs68L_reg[5][5] (.clk (\Clks[clk] ), .d (n_5336), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [5]));
  CDN_flop \regs68L_reg[5][6] (.clk (\Clks[clk] ), .d (n_5337), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [6]));
  CDN_flop \regs68L_reg[5][7] (.clk (\Clks[clk] ), .d (n_5338), .sena
       (n_5331), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [7]));
  CDN_flop \regs68L_reg[5][8] (.clk (\Clks[clk] ), .d (n_5339), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [8]));
  CDN_flop \regs68L_reg[5][9] (.clk (\Clks[clk] ), .d (n_5341), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [9]));
  CDN_flop \regs68L_reg[5][10] (.clk (\Clks[clk] ), .d (n_5342), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [10]));
  CDN_flop \regs68L_reg[5][11] (.clk (\Clks[clk] ), .d (n_5343), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [11]));
  CDN_flop \regs68L_reg[5][12] (.clk (\Clks[clk] ), .d (n_5344), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [12]));
  CDN_flop \regs68L_reg[5][13] (.clk (\Clks[clk] ), .d (n_5345), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [13]));
  CDN_flop \regs68L_reg[5][14] (.clk (\Clks[clk] ), .d (n_5346), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [14]));
  CDN_flop \regs68L_reg[5][15] (.clk (\Clks[clk] ), .d (n_5347), .sena
       (n_5340), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[5] [15]));
  CDN_flop \regs68L_reg[4][0] (.clk (\Clks[clk] ), .d (n_5409), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [0]));
  CDN_flop \regs68L_reg[4][1] (.clk (\Clks[clk] ), .d (n_5411), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [1]));
  CDN_flop \regs68L_reg[4][2] (.clk (\Clks[clk] ), .d (n_5412), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [2]));
  CDN_flop \regs68L_reg[4][3] (.clk (\Clks[clk] ), .d (n_5413), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [3]));
  CDN_flop \regs68L_reg[4][4] (.clk (\Clks[clk] ), .d (n_5414), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [4]));
  CDN_flop \regs68L_reg[4][5] (.clk (\Clks[clk] ), .d (n_5415), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [5]));
  CDN_flop \regs68L_reg[4][6] (.clk (\Clks[clk] ), .d (n_5416), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [6]));
  CDN_flop \regs68L_reg[4][7] (.clk (\Clks[clk] ), .d (n_5417), .sena
       (n_5410), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [7]));
  CDN_flop \regs68L_reg[4][8] (.clk (\Clks[clk] ), .d (n_5418), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [8]));
  CDN_flop \regs68L_reg[4][9] (.clk (\Clks[clk] ), .d (n_5420), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [9]));
  CDN_flop \regs68L_reg[4][10] (.clk (\Clks[clk] ), .d (n_5421), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [10]));
  CDN_flop \regs68L_reg[4][11] (.clk (\Clks[clk] ), .d (n_5422), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [11]));
  CDN_flop \regs68L_reg[4][12] (.clk (\Clks[clk] ), .d (n_5423), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [12]));
  CDN_flop \regs68L_reg[4][13] (.clk (\Clks[clk] ), .d (n_5424), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [13]));
  CDN_flop \regs68L_reg[4][14] (.clk (\Clks[clk] ), .d (n_5425), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [14]));
  CDN_flop \regs68L_reg[4][15] (.clk (\Clks[clk] ), .d (n_5426), .sena
       (n_5419), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[4] [15]));
  CDN_flop \regs68L_reg[3][0] (.clk (\Clks[clk] ), .d (n_5488), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [0]));
  CDN_flop \regs68L_reg[3][1] (.clk (\Clks[clk] ), .d (n_5490), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [1]));
  CDN_flop \regs68L_reg[3][2] (.clk (\Clks[clk] ), .d (n_5491), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [2]));
  CDN_flop \regs68L_reg[3][3] (.clk (\Clks[clk] ), .d (n_5492), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [3]));
  CDN_flop \regs68L_reg[3][4] (.clk (\Clks[clk] ), .d (n_5493), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [4]));
  CDN_flop \regs68L_reg[3][5] (.clk (\Clks[clk] ), .d (n_5494), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [5]));
  CDN_flop \regs68L_reg[3][6] (.clk (\Clks[clk] ), .d (n_5495), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [6]));
  CDN_flop \regs68L_reg[3][7] (.clk (\Clks[clk] ), .d (n_5496), .sena
       (n_5489), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [7]));
  CDN_flop \regs68L_reg[3][8] (.clk (\Clks[clk] ), .d (n_5497), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [8]));
  CDN_flop \regs68L_reg[3][9] (.clk (\Clks[clk] ), .d (n_5499), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [9]));
  CDN_flop \regs68L_reg[3][10] (.clk (\Clks[clk] ), .d (n_5500), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [10]));
  CDN_flop \regs68L_reg[3][11] (.clk (\Clks[clk] ), .d (n_5501), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [11]));
  CDN_flop \regs68L_reg[3][12] (.clk (\Clks[clk] ), .d (n_5502), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [12]));
  CDN_flop \regs68L_reg[3][13] (.clk (\Clks[clk] ), .d (n_5503), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [13]));
  CDN_flop \regs68L_reg[3][14] (.clk (\Clks[clk] ), .d (n_5504), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [14]));
  CDN_flop \regs68L_reg[3][15] (.clk (\Clks[clk] ), .d (n_5505), .sena
       (n_5498), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[3] [15]));
  CDN_flop \regs68L_reg[2][0] (.clk (\Clks[clk] ), .d (n_5567), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [0]));
  CDN_flop \regs68L_reg[2][1] (.clk (\Clks[clk] ), .d (n_5569), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [1]));
  CDN_flop \regs68L_reg[2][2] (.clk (\Clks[clk] ), .d (n_5570), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [2]));
  CDN_flop \regs68L_reg[2][3] (.clk (\Clks[clk] ), .d (n_5571), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [3]));
  CDN_flop \regs68L_reg[2][4] (.clk (\Clks[clk] ), .d (n_5572), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [4]));
  CDN_flop \regs68L_reg[2][5] (.clk (\Clks[clk] ), .d (n_5573), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [5]));
  CDN_flop \regs68L_reg[2][6] (.clk (\Clks[clk] ), .d (n_5574), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [6]));
  CDN_flop \regs68L_reg[2][7] (.clk (\Clks[clk] ), .d (n_5575), .sena
       (n_5568), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [7]));
  CDN_flop \regs68L_reg[2][8] (.clk (\Clks[clk] ), .d (n_5576), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [8]));
  CDN_flop \regs68L_reg[2][9] (.clk (\Clks[clk] ), .d (n_5578), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [9]));
  CDN_flop \regs68L_reg[2][10] (.clk (\Clks[clk] ), .d (n_5579), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [10]));
  CDN_flop \regs68L_reg[2][11] (.clk (\Clks[clk] ), .d (n_5580), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [11]));
  CDN_flop \regs68L_reg[2][12] (.clk (\Clks[clk] ), .d (n_5581), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [12]));
  CDN_flop \regs68L_reg[2][13] (.clk (\Clks[clk] ), .d (n_5582), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [13]));
  CDN_flop \regs68L_reg[2][14] (.clk (\Clks[clk] ), .d (n_5583), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [14]));
  CDN_flop \regs68L_reg[2][15] (.clk (\Clks[clk] ), .d (n_5584), .sena
       (n_5577), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[2] [15]));
  CDN_flop \regs68L_reg[1][0] (.clk (\Clks[clk] ), .d (n_5646), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [0]));
  CDN_flop \regs68L_reg[1][1] (.clk (\Clks[clk] ), .d (n_5648), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [1]));
  CDN_flop \regs68L_reg[1][2] (.clk (\Clks[clk] ), .d (n_5649), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [2]));
  CDN_flop \regs68L_reg[1][3] (.clk (\Clks[clk] ), .d (n_5650), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [3]));
  CDN_flop \regs68L_reg[1][4] (.clk (\Clks[clk] ), .d (n_5651), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [4]));
  CDN_flop \regs68L_reg[1][5] (.clk (\Clks[clk] ), .d (n_5652), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [5]));
  CDN_flop \regs68L_reg[1][6] (.clk (\Clks[clk] ), .d (n_5653), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [6]));
  CDN_flop \regs68L_reg[1][7] (.clk (\Clks[clk] ), .d (n_5654), .sena
       (n_5647), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [7]));
  CDN_flop \regs68L_reg[1][8] (.clk (\Clks[clk] ), .d (n_5655), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [8]));
  CDN_flop \regs68L_reg[1][9] (.clk (\Clks[clk] ), .d (n_5657), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [9]));
  CDN_flop \regs68L_reg[1][10] (.clk (\Clks[clk] ), .d (n_5658), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [10]));
  CDN_flop \regs68L_reg[1][11] (.clk (\Clks[clk] ), .d (n_5659), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [11]));
  CDN_flop \regs68L_reg[1][12] (.clk (\Clks[clk] ), .d (n_5660), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [12]));
  CDN_flop \regs68L_reg[1][13] (.clk (\Clks[clk] ), .d (n_5661), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [13]));
  CDN_flop \regs68L_reg[1][14] (.clk (\Clks[clk] ), .d (n_5662), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [14]));
  CDN_flop \regs68L_reg[1][15] (.clk (\Clks[clk] ), .d (n_5663), .sena
       (n_5656), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[1] [15]));
  CDN_flop \regs68L_reg[0][0] (.clk (\Clks[clk] ), .d (n_5725), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [0]));
  CDN_flop \regs68L_reg[0][1] (.clk (\Clks[clk] ), .d (n_5727), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [1]));
  CDN_flop \regs68L_reg[0][2] (.clk (\Clks[clk] ), .d (n_5728), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [2]));
  CDN_flop \regs68L_reg[0][3] (.clk (\Clks[clk] ), .d (n_5729), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [3]));
  CDN_flop \regs68L_reg[0][4] (.clk (\Clks[clk] ), .d (n_5730), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [4]));
  CDN_flop \regs68L_reg[0][5] (.clk (\Clks[clk] ), .d (n_5731), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [5]));
  CDN_flop \regs68L_reg[0][6] (.clk (\Clks[clk] ), .d (n_5732), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [6]));
  CDN_flop \regs68L_reg[0][7] (.clk (\Clks[clk] ), .d (n_5733), .sena
       (n_5726), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [7]));
  CDN_flop \regs68L_reg[0][8] (.clk (\Clks[clk] ), .d (n_5734), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [8]));
  CDN_flop \regs68L_reg[0][9] (.clk (\Clks[clk] ), .d (n_5736), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [9]));
  CDN_flop \regs68L_reg[0][10] (.clk (\Clks[clk] ), .d (n_5737), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [10]));
  CDN_flop \regs68L_reg[0][11] (.clk (\Clks[clk] ), .d (n_5738), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [11]));
  CDN_flop \regs68L_reg[0][12] (.clk (\Clks[clk] ), .d (n_5739), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [12]));
  CDN_flop \regs68L_reg[0][13] (.clk (\Clks[clk] ), .d (n_5740), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [13]));
  CDN_flop \regs68L_reg[0][14] (.clk (\Clks[clk] ), .d (n_5741), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [14]));
  CDN_flop \regs68L_reg[0][15] (.clk (\Clks[clk] ), .d (n_5742), .sena
       (n_5735), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68L[0] [15]));
  CDN_flop \regs68H_reg[17][0] (.clk (\Clks[clk] ), .d (n_5751), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [0]));
  CDN_flop \regs68H_reg[17][1] (.clk (\Clks[clk] ), .d (n_5753), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [1]));
  CDN_flop \regs68H_reg[17][2] (.clk (\Clks[clk] ), .d (n_5754), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [2]));
  CDN_flop \regs68H_reg[17][3] (.clk (\Clks[clk] ), .d (n_5755), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [3]));
  CDN_flop \regs68H_reg[17][4] (.clk (\Clks[clk] ), .d (n_5756), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [4]));
  CDN_flop \regs68H_reg[17][5] (.clk (\Clks[clk] ), .d (n_5757), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [5]));
  CDN_flop \regs68H_reg[17][6] (.clk (\Clks[clk] ), .d (n_5758), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [6]));
  CDN_flop \regs68H_reg[17][7] (.clk (\Clks[clk] ), .d (n_5759), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [7]));
  CDN_flop \regs68H_reg[17][8] (.clk (\Clks[clk] ), .d (n_5760), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [8]));
  CDN_flop \regs68H_reg[17][9] (.clk (\Clks[clk] ), .d (n_5761), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [9]));
  CDN_flop \regs68H_reg[17][10] (.clk (\Clks[clk] ), .d (n_5762), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [10]));
  CDN_flop \regs68H_reg[17][11] (.clk (\Clks[clk] ), .d (n_5763), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [11]));
  CDN_flop \regs68H_reg[17][12] (.clk (\Clks[clk] ), .d (n_5764), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [12]));
  CDN_flop \regs68H_reg[17][13] (.clk (\Clks[clk] ), .d (n_5765), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [13]));
  CDN_flop \regs68H_reg[17][14] (.clk (\Clks[clk] ), .d (n_5766), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [14]));
  CDN_flop \regs68H_reg[17][15] (.clk (\Clks[clk] ), .d (n_5767), .sena
       (n_5752), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[17] [15]));
  CDN_flop \regs68H_reg[16][0] (.clk (\Clks[clk] ), .d (n_5775), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [0]));
  CDN_flop \regs68H_reg[16][1] (.clk (\Clks[clk] ), .d (n_5777), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [1]));
  CDN_flop \regs68H_reg[16][2] (.clk (\Clks[clk] ), .d (n_5778), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [2]));
  CDN_flop \regs68H_reg[16][3] (.clk (\Clks[clk] ), .d (n_5779), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [3]));
  CDN_flop \regs68H_reg[16][4] (.clk (\Clks[clk] ), .d (n_5780), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [4]));
  CDN_flop \regs68H_reg[16][5] (.clk (\Clks[clk] ), .d (n_5781), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [5]));
  CDN_flop \regs68H_reg[16][6] (.clk (\Clks[clk] ), .d (n_5782), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [6]));
  CDN_flop \regs68H_reg[16][7] (.clk (\Clks[clk] ), .d (n_5783), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [7]));
  CDN_flop \regs68H_reg[16][8] (.clk (\Clks[clk] ), .d (n_5784), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [8]));
  CDN_flop \regs68H_reg[16][9] (.clk (\Clks[clk] ), .d (n_5785), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [9]));
  CDN_flop \regs68H_reg[16][10] (.clk (\Clks[clk] ), .d (n_5786), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [10]));
  CDN_flop \regs68H_reg[16][11] (.clk (\Clks[clk] ), .d (n_5787), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [11]));
  CDN_flop \regs68H_reg[16][12] (.clk (\Clks[clk] ), .d (n_5788), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [12]));
  CDN_flop \regs68H_reg[16][13] (.clk (\Clks[clk] ), .d (n_5789), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [13]));
  CDN_flop \regs68H_reg[16][14] (.clk (\Clks[clk] ), .d (n_5790), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [14]));
  CDN_flop \regs68H_reg[16][15] (.clk (\Clks[clk] ), .d (n_5791), .sena
       (n_5776), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[16] [15]));
  CDN_flop \regs68H_reg[15][0] (.clk (\Clks[clk] ), .d (n_5799), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [0]));
  CDN_flop \regs68H_reg[15][1] (.clk (\Clks[clk] ), .d (n_5801), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [1]));
  CDN_flop \regs68H_reg[15][2] (.clk (\Clks[clk] ), .d (n_5802), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [2]));
  CDN_flop \regs68H_reg[15][3] (.clk (\Clks[clk] ), .d (n_5803), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [3]));
  CDN_flop \regs68H_reg[15][4] (.clk (\Clks[clk] ), .d (n_5804), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [4]));
  CDN_flop \regs68H_reg[15][5] (.clk (\Clks[clk] ), .d (n_5805), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [5]));
  CDN_flop \regs68H_reg[15][6] (.clk (\Clks[clk] ), .d (n_5806), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [6]));
  CDN_flop \regs68H_reg[15][7] (.clk (\Clks[clk] ), .d (n_5807), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [7]));
  CDN_flop \regs68H_reg[15][8] (.clk (\Clks[clk] ), .d (n_5808), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [8]));
  CDN_flop \regs68H_reg[15][9] (.clk (\Clks[clk] ), .d (n_5809), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [9]));
  CDN_flop \regs68H_reg[15][10] (.clk (\Clks[clk] ), .d (n_5810), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [10]));
  CDN_flop \regs68H_reg[15][11] (.clk (\Clks[clk] ), .d (n_5811), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [11]));
  CDN_flop \regs68H_reg[15][12] (.clk (\Clks[clk] ), .d (n_5812), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [12]));
  CDN_flop \regs68H_reg[15][13] (.clk (\Clks[clk] ), .d (n_5813), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [13]));
  CDN_flop \regs68H_reg[15][14] (.clk (\Clks[clk] ), .d (n_5814), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [14]));
  CDN_flop \regs68H_reg[15][15] (.clk (\Clks[clk] ), .d (n_5815), .sena
       (n_5800), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[15] [15]));
  CDN_flop \regs68H_reg[14][0] (.clk (\Clks[clk] ), .d (n_5823), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [0]));
  CDN_flop \regs68H_reg[14][1] (.clk (\Clks[clk] ), .d (n_5825), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [1]));
  CDN_flop \regs68H_reg[14][2] (.clk (\Clks[clk] ), .d (n_5826), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [2]));
  CDN_flop \regs68H_reg[14][3] (.clk (\Clks[clk] ), .d (n_5827), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [3]));
  CDN_flop \regs68H_reg[14][4] (.clk (\Clks[clk] ), .d (n_5828), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [4]));
  CDN_flop \regs68H_reg[14][5] (.clk (\Clks[clk] ), .d (n_5829), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [5]));
  CDN_flop \regs68H_reg[14][6] (.clk (\Clks[clk] ), .d (n_5830), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [6]));
  CDN_flop \regs68H_reg[14][7] (.clk (\Clks[clk] ), .d (n_5831), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [7]));
  CDN_flop \regs68H_reg[14][8] (.clk (\Clks[clk] ), .d (n_5832), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [8]));
  CDN_flop \regs68H_reg[14][9] (.clk (\Clks[clk] ), .d (n_5833), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [9]));
  CDN_flop \regs68H_reg[14][10] (.clk (\Clks[clk] ), .d (n_5834), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [10]));
  CDN_flop \regs68H_reg[14][11] (.clk (\Clks[clk] ), .d (n_5835), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [11]));
  CDN_flop \regs68H_reg[14][12] (.clk (\Clks[clk] ), .d (n_5836), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [12]));
  CDN_flop \regs68H_reg[14][13] (.clk (\Clks[clk] ), .d (n_5837), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [13]));
  CDN_flop \regs68H_reg[14][14] (.clk (\Clks[clk] ), .d (n_5838), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [14]));
  CDN_flop \regs68H_reg[14][15] (.clk (\Clks[clk] ), .d (n_5839), .sena
       (n_5824), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[14] [15]));
  CDN_flop \regs68H_reg[13][0] (.clk (\Clks[clk] ), .d (n_5847), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [0]));
  CDN_flop \regs68H_reg[13][1] (.clk (\Clks[clk] ), .d (n_5849), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [1]));
  CDN_flop \regs68H_reg[13][2] (.clk (\Clks[clk] ), .d (n_5850), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [2]));
  CDN_flop \regs68H_reg[13][3] (.clk (\Clks[clk] ), .d (n_5851), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [3]));
  CDN_flop \regs68H_reg[13][4] (.clk (\Clks[clk] ), .d (n_5852), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [4]));
  CDN_flop \regs68H_reg[13][5] (.clk (\Clks[clk] ), .d (n_5853), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [5]));
  CDN_flop \regs68H_reg[13][6] (.clk (\Clks[clk] ), .d (n_5854), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [6]));
  CDN_flop \regs68H_reg[13][7] (.clk (\Clks[clk] ), .d (n_5855), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [7]));
  CDN_flop \regs68H_reg[13][8] (.clk (\Clks[clk] ), .d (n_5856), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [8]));
  CDN_flop \regs68H_reg[13][9] (.clk (\Clks[clk] ), .d (n_5857), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [9]));
  CDN_flop \regs68H_reg[13][10] (.clk (\Clks[clk] ), .d (n_5858), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [10]));
  CDN_flop \regs68H_reg[13][11] (.clk (\Clks[clk] ), .d (n_5859), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [11]));
  CDN_flop \regs68H_reg[13][12] (.clk (\Clks[clk] ), .d (n_5860), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [12]));
  CDN_flop \regs68H_reg[13][13] (.clk (\Clks[clk] ), .d (n_5861), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [13]));
  CDN_flop \regs68H_reg[13][14] (.clk (\Clks[clk] ), .d (n_5862), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [14]));
  CDN_flop \regs68H_reg[13][15] (.clk (\Clks[clk] ), .d (n_5863), .sena
       (n_5848), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[13] [15]));
  CDN_flop \regs68H_reg[12][0] (.clk (\Clks[clk] ), .d (n_5871), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [0]));
  CDN_flop \regs68H_reg[12][1] (.clk (\Clks[clk] ), .d (n_5873), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [1]));
  CDN_flop \regs68H_reg[12][2] (.clk (\Clks[clk] ), .d (n_5874), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [2]));
  CDN_flop \regs68H_reg[12][3] (.clk (\Clks[clk] ), .d (n_5875), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [3]));
  CDN_flop \regs68H_reg[12][4] (.clk (\Clks[clk] ), .d (n_5876), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [4]));
  CDN_flop \regs68H_reg[12][5] (.clk (\Clks[clk] ), .d (n_5877), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [5]));
  CDN_flop \regs68H_reg[12][6] (.clk (\Clks[clk] ), .d (n_5878), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [6]));
  CDN_flop \regs68H_reg[12][7] (.clk (\Clks[clk] ), .d (n_5879), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [7]));
  CDN_flop \regs68H_reg[12][8] (.clk (\Clks[clk] ), .d (n_5880), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [8]));
  CDN_flop \regs68H_reg[12][9] (.clk (\Clks[clk] ), .d (n_5881), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [9]));
  CDN_flop \regs68H_reg[12][10] (.clk (\Clks[clk] ), .d (n_5882), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [10]));
  CDN_flop \regs68H_reg[12][11] (.clk (\Clks[clk] ), .d (n_5883), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [11]));
  CDN_flop \regs68H_reg[12][12] (.clk (\Clks[clk] ), .d (n_5884), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [12]));
  CDN_flop \regs68H_reg[12][13] (.clk (\Clks[clk] ), .d (n_5885), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [13]));
  CDN_flop \regs68H_reg[12][14] (.clk (\Clks[clk] ), .d (n_5886), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [14]));
  CDN_flop \regs68H_reg[12][15] (.clk (\Clks[clk] ), .d (n_5887), .sena
       (n_5872), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[12] [15]));
  CDN_flop \regs68H_reg[11][0] (.clk (\Clks[clk] ), .d (n_5895), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [0]));
  CDN_flop \regs68H_reg[11][1] (.clk (\Clks[clk] ), .d (n_5897), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [1]));
  CDN_flop \regs68H_reg[11][2] (.clk (\Clks[clk] ), .d (n_5898), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [2]));
  CDN_flop \regs68H_reg[11][3] (.clk (\Clks[clk] ), .d (n_5899), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [3]));
  CDN_flop \regs68H_reg[11][4] (.clk (\Clks[clk] ), .d (n_5900), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [4]));
  CDN_flop \regs68H_reg[11][5] (.clk (\Clks[clk] ), .d (n_5901), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [5]));
  CDN_flop \regs68H_reg[11][6] (.clk (\Clks[clk] ), .d (n_5902), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [6]));
  CDN_flop \regs68H_reg[11][7] (.clk (\Clks[clk] ), .d (n_5903), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [7]));
  CDN_flop \regs68H_reg[11][8] (.clk (\Clks[clk] ), .d (n_5904), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [8]));
  CDN_flop \regs68H_reg[11][9] (.clk (\Clks[clk] ), .d (n_5905), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [9]));
  CDN_flop \regs68H_reg[11][10] (.clk (\Clks[clk] ), .d (n_5906), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [10]));
  CDN_flop \regs68H_reg[11][11] (.clk (\Clks[clk] ), .d (n_5907), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [11]));
  CDN_flop \regs68H_reg[11][12] (.clk (\Clks[clk] ), .d (n_5908), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [12]));
  CDN_flop \regs68H_reg[11][13] (.clk (\Clks[clk] ), .d (n_5909), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [13]));
  CDN_flop \regs68H_reg[11][14] (.clk (\Clks[clk] ), .d (n_5910), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [14]));
  CDN_flop \regs68H_reg[11][15] (.clk (\Clks[clk] ), .d (n_5911), .sena
       (n_5896), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[11] [15]));
  CDN_flop \regs68H_reg[10][0] (.clk (\Clks[clk] ), .d (n_5919), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [0]));
  CDN_flop \regs68H_reg[10][1] (.clk (\Clks[clk] ), .d (n_5921), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [1]));
  CDN_flop \regs68H_reg[10][2] (.clk (\Clks[clk] ), .d (n_5922), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [2]));
  CDN_flop \regs68H_reg[10][3] (.clk (\Clks[clk] ), .d (n_5923), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [3]));
  CDN_flop \regs68H_reg[10][4] (.clk (\Clks[clk] ), .d (n_5924), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [4]));
  CDN_flop \regs68H_reg[10][5] (.clk (\Clks[clk] ), .d (n_5925), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [5]));
  CDN_flop \regs68H_reg[10][6] (.clk (\Clks[clk] ), .d (n_5926), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [6]));
  CDN_flop \regs68H_reg[10][7] (.clk (\Clks[clk] ), .d (n_5927), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [7]));
  CDN_flop \regs68H_reg[10][8] (.clk (\Clks[clk] ), .d (n_5928), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [8]));
  CDN_flop \regs68H_reg[10][9] (.clk (\Clks[clk] ), .d (n_5929), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [9]));
  CDN_flop \regs68H_reg[10][10] (.clk (\Clks[clk] ), .d (n_5930), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [10]));
  CDN_flop \regs68H_reg[10][11] (.clk (\Clks[clk] ), .d (n_5931), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [11]));
  CDN_flop \regs68H_reg[10][12] (.clk (\Clks[clk] ), .d (n_5932), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [12]));
  CDN_flop \regs68H_reg[10][13] (.clk (\Clks[clk] ), .d (n_5933), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [13]));
  CDN_flop \regs68H_reg[10][14] (.clk (\Clks[clk] ), .d (n_5934), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [14]));
  CDN_flop \regs68H_reg[10][15] (.clk (\Clks[clk] ), .d (n_5935), .sena
       (n_5920), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[10] [15]));
  CDN_flop \regs68H_reg[9][0] (.clk (\Clks[clk] ), .d (n_5943), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [0]));
  CDN_flop \regs68H_reg[9][1] (.clk (\Clks[clk] ), .d (n_5945), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [1]));
  CDN_flop \regs68H_reg[9][2] (.clk (\Clks[clk] ), .d (n_5946), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [2]));
  CDN_flop \regs68H_reg[9][3] (.clk (\Clks[clk] ), .d (n_5947), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [3]));
  CDN_flop \regs68H_reg[9][4] (.clk (\Clks[clk] ), .d (n_5948), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [4]));
  CDN_flop \regs68H_reg[9][5] (.clk (\Clks[clk] ), .d (n_5949), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [5]));
  CDN_flop \regs68H_reg[9][6] (.clk (\Clks[clk] ), .d (n_5950), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [6]));
  CDN_flop \regs68H_reg[9][7] (.clk (\Clks[clk] ), .d (n_5951), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [7]));
  CDN_flop \regs68H_reg[9][8] (.clk (\Clks[clk] ), .d (n_5952), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [8]));
  CDN_flop \regs68H_reg[9][9] (.clk (\Clks[clk] ), .d (n_5953), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [9]));
  CDN_flop \regs68H_reg[9][10] (.clk (\Clks[clk] ), .d (n_5954), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [10]));
  CDN_flop \regs68H_reg[9][11] (.clk (\Clks[clk] ), .d (n_5955), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [11]));
  CDN_flop \regs68H_reg[9][12] (.clk (\Clks[clk] ), .d (n_5956), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [12]));
  CDN_flop \regs68H_reg[9][13] (.clk (\Clks[clk] ), .d (n_5957), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [13]));
  CDN_flop \regs68H_reg[9][14] (.clk (\Clks[clk] ), .d (n_5958), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [14]));
  CDN_flop \regs68H_reg[9][15] (.clk (\Clks[clk] ), .d (n_5959), .sena
       (n_5944), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[9] [15]));
  CDN_flop \regs68H_reg[8][0] (.clk (\Clks[clk] ), .d (n_5967), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [0]));
  CDN_flop \regs68H_reg[8][1] (.clk (\Clks[clk] ), .d (n_5969), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [1]));
  CDN_flop \regs68H_reg[8][2] (.clk (\Clks[clk] ), .d (n_5970), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [2]));
  CDN_flop \regs68H_reg[8][3] (.clk (\Clks[clk] ), .d (n_5971), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [3]));
  CDN_flop \regs68H_reg[8][4] (.clk (\Clks[clk] ), .d (n_5972), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [4]));
  CDN_flop \regs68H_reg[8][5] (.clk (\Clks[clk] ), .d (n_5973), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [5]));
  CDN_flop \regs68H_reg[8][6] (.clk (\Clks[clk] ), .d (n_5974), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [6]));
  CDN_flop \regs68H_reg[8][7] (.clk (\Clks[clk] ), .d (n_5975), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [7]));
  CDN_flop \regs68H_reg[8][8] (.clk (\Clks[clk] ), .d (n_5976), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [8]));
  CDN_flop \regs68H_reg[8][9] (.clk (\Clks[clk] ), .d (n_5977), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [9]));
  CDN_flop \regs68H_reg[8][10] (.clk (\Clks[clk] ), .d (n_5978), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [10]));
  CDN_flop \regs68H_reg[8][11] (.clk (\Clks[clk] ), .d (n_5979), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [11]));
  CDN_flop \regs68H_reg[8][12] (.clk (\Clks[clk] ), .d (n_5980), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [12]));
  CDN_flop \regs68H_reg[8][13] (.clk (\Clks[clk] ), .d (n_5981), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [13]));
  CDN_flop \regs68H_reg[8][14] (.clk (\Clks[clk] ), .d (n_5982), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [14]));
  CDN_flop \regs68H_reg[8][15] (.clk (\Clks[clk] ), .d (n_5983), .sena
       (n_5968), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[8] [15]));
  CDN_flop \regs68H_reg[7][0] (.clk (\Clks[clk] ), .d (n_5991), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [0]));
  CDN_flop \regs68H_reg[7][1] (.clk (\Clks[clk] ), .d (n_5993), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [1]));
  CDN_flop \regs68H_reg[7][2] (.clk (\Clks[clk] ), .d (n_5994), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [2]));
  CDN_flop \regs68H_reg[7][3] (.clk (\Clks[clk] ), .d (n_5995), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [3]));
  CDN_flop \regs68H_reg[7][4] (.clk (\Clks[clk] ), .d (n_5996), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [4]));
  CDN_flop \regs68H_reg[7][5] (.clk (\Clks[clk] ), .d (n_5997), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [5]));
  CDN_flop \regs68H_reg[7][6] (.clk (\Clks[clk] ), .d (n_5998), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [6]));
  CDN_flop \regs68H_reg[7][7] (.clk (\Clks[clk] ), .d (n_5999), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [7]));
  CDN_flop \regs68H_reg[7][8] (.clk (\Clks[clk] ), .d (n_6000), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [8]));
  CDN_flop \regs68H_reg[7][9] (.clk (\Clks[clk] ), .d (n_6001), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [9]));
  CDN_flop \regs68H_reg[7][10] (.clk (\Clks[clk] ), .d (n_6002), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [10]));
  CDN_flop \regs68H_reg[7][11] (.clk (\Clks[clk] ), .d (n_6003), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [11]));
  CDN_flop \regs68H_reg[7][12] (.clk (\Clks[clk] ), .d (n_6004), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [12]));
  CDN_flop \regs68H_reg[7][13] (.clk (\Clks[clk] ), .d (n_6005), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [13]));
  CDN_flop \regs68H_reg[7][14] (.clk (\Clks[clk] ), .d (n_6006), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [14]));
  CDN_flop \regs68H_reg[7][15] (.clk (\Clks[clk] ), .d (n_6007), .sena
       (n_5992), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[7] [15]));
  CDN_flop \regs68H_reg[6][0] (.clk (\Clks[clk] ), .d (n_6015), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [0]));
  CDN_flop \regs68H_reg[6][1] (.clk (\Clks[clk] ), .d (n_6017), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [1]));
  CDN_flop \regs68H_reg[6][2] (.clk (\Clks[clk] ), .d (n_6018), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [2]));
  CDN_flop \regs68H_reg[6][3] (.clk (\Clks[clk] ), .d (n_6019), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [3]));
  CDN_flop \regs68H_reg[6][4] (.clk (\Clks[clk] ), .d (n_6020), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [4]));
  CDN_flop \regs68H_reg[6][5] (.clk (\Clks[clk] ), .d (n_6021), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [5]));
  CDN_flop \regs68H_reg[6][6] (.clk (\Clks[clk] ), .d (n_6022), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [6]));
  CDN_flop \regs68H_reg[6][7] (.clk (\Clks[clk] ), .d (n_6023), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [7]));
  CDN_flop \regs68H_reg[6][8] (.clk (\Clks[clk] ), .d (n_6024), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [8]));
  CDN_flop \regs68H_reg[6][9] (.clk (\Clks[clk] ), .d (n_6025), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [9]));
  CDN_flop \regs68H_reg[6][10] (.clk (\Clks[clk] ), .d (n_6026), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [10]));
  CDN_flop \regs68H_reg[6][11] (.clk (\Clks[clk] ), .d (n_6027), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [11]));
  CDN_flop \regs68H_reg[6][12] (.clk (\Clks[clk] ), .d (n_6028), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [12]));
  CDN_flop \regs68H_reg[6][13] (.clk (\Clks[clk] ), .d (n_6029), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [13]));
  CDN_flop \regs68H_reg[6][14] (.clk (\Clks[clk] ), .d (n_6030), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [14]));
  CDN_flop \regs68H_reg[6][15] (.clk (\Clks[clk] ), .d (n_6031), .sena
       (n_6016), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[6] [15]));
  CDN_flop \regs68H_reg[5][0] (.clk (\Clks[clk] ), .d (n_6039), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [0]));
  CDN_flop \regs68H_reg[5][1] (.clk (\Clks[clk] ), .d (n_6041), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [1]));
  CDN_flop \regs68H_reg[5][2] (.clk (\Clks[clk] ), .d (n_6042), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [2]));
  CDN_flop \regs68H_reg[5][3] (.clk (\Clks[clk] ), .d (n_6043), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [3]));
  CDN_flop \regs68H_reg[5][4] (.clk (\Clks[clk] ), .d (n_6044), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [4]));
  CDN_flop \regs68H_reg[5][5] (.clk (\Clks[clk] ), .d (n_6045), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [5]));
  CDN_flop \regs68H_reg[5][6] (.clk (\Clks[clk] ), .d (n_6046), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [6]));
  CDN_flop \regs68H_reg[5][7] (.clk (\Clks[clk] ), .d (n_6047), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [7]));
  CDN_flop \regs68H_reg[5][8] (.clk (\Clks[clk] ), .d (n_6048), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [8]));
  CDN_flop \regs68H_reg[5][9] (.clk (\Clks[clk] ), .d (n_6049), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [9]));
  CDN_flop \regs68H_reg[5][10] (.clk (\Clks[clk] ), .d (n_6050), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [10]));
  CDN_flop \regs68H_reg[5][11] (.clk (\Clks[clk] ), .d (n_6051), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [11]));
  CDN_flop \regs68H_reg[5][12] (.clk (\Clks[clk] ), .d (n_6052), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [12]));
  CDN_flop \regs68H_reg[5][13] (.clk (\Clks[clk] ), .d (n_6053), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [13]));
  CDN_flop \regs68H_reg[5][14] (.clk (\Clks[clk] ), .d (n_6054), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [14]));
  CDN_flop \regs68H_reg[5][15] (.clk (\Clks[clk] ), .d (n_6055), .sena
       (n_6040), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[5] [15]));
  CDN_flop \regs68H_reg[4][0] (.clk (\Clks[clk] ), .d (n_6063), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [0]));
  CDN_flop \regs68H_reg[4][1] (.clk (\Clks[clk] ), .d (n_6065), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [1]));
  CDN_flop \regs68H_reg[4][2] (.clk (\Clks[clk] ), .d (n_6066), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [2]));
  CDN_flop \regs68H_reg[4][3] (.clk (\Clks[clk] ), .d (n_6067), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [3]));
  CDN_flop \regs68H_reg[4][4] (.clk (\Clks[clk] ), .d (n_6068), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [4]));
  CDN_flop \regs68H_reg[4][5] (.clk (\Clks[clk] ), .d (n_6069), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [5]));
  CDN_flop \regs68H_reg[4][6] (.clk (\Clks[clk] ), .d (n_6070), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [6]));
  CDN_flop \regs68H_reg[4][7] (.clk (\Clks[clk] ), .d (n_6071), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [7]));
  CDN_flop \regs68H_reg[4][8] (.clk (\Clks[clk] ), .d (n_6072), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [8]));
  CDN_flop \regs68H_reg[4][9] (.clk (\Clks[clk] ), .d (n_6073), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [9]));
  CDN_flop \regs68H_reg[4][10] (.clk (\Clks[clk] ), .d (n_6074), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [10]));
  CDN_flop \regs68H_reg[4][11] (.clk (\Clks[clk] ), .d (n_6075), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [11]));
  CDN_flop \regs68H_reg[4][12] (.clk (\Clks[clk] ), .d (n_6076), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [12]));
  CDN_flop \regs68H_reg[4][13] (.clk (\Clks[clk] ), .d (n_6077), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [13]));
  CDN_flop \regs68H_reg[4][14] (.clk (\Clks[clk] ), .d (n_6078), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [14]));
  CDN_flop \regs68H_reg[4][15] (.clk (\Clks[clk] ), .d (n_6079), .sena
       (n_6064), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[4] [15]));
  CDN_flop \regs68H_reg[3][0] (.clk (\Clks[clk] ), .d (n_6087), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [0]));
  CDN_flop \regs68H_reg[3][1] (.clk (\Clks[clk] ), .d (n_6089), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [1]));
  CDN_flop \regs68H_reg[3][2] (.clk (\Clks[clk] ), .d (n_6090), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [2]));
  CDN_flop \regs68H_reg[3][3] (.clk (\Clks[clk] ), .d (n_6091), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [3]));
  CDN_flop \regs68H_reg[3][4] (.clk (\Clks[clk] ), .d (n_6092), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [4]));
  CDN_flop \regs68H_reg[3][5] (.clk (\Clks[clk] ), .d (n_6093), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [5]));
  CDN_flop \regs68H_reg[3][6] (.clk (\Clks[clk] ), .d (n_6094), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [6]));
  CDN_flop \regs68H_reg[3][7] (.clk (\Clks[clk] ), .d (n_6095), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [7]));
  CDN_flop \regs68H_reg[3][8] (.clk (\Clks[clk] ), .d (n_6096), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [8]));
  CDN_flop \regs68H_reg[3][9] (.clk (\Clks[clk] ), .d (n_6097), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [9]));
  CDN_flop \regs68H_reg[3][10] (.clk (\Clks[clk] ), .d (n_6098), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [10]));
  CDN_flop \regs68H_reg[3][11] (.clk (\Clks[clk] ), .d (n_6099), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [11]));
  CDN_flop \regs68H_reg[3][12] (.clk (\Clks[clk] ), .d (n_6100), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [12]));
  CDN_flop \regs68H_reg[3][13] (.clk (\Clks[clk] ), .d (n_6101), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [13]));
  CDN_flop \regs68H_reg[3][14] (.clk (\Clks[clk] ), .d (n_6102), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [14]));
  CDN_flop \regs68H_reg[3][15] (.clk (\Clks[clk] ), .d (n_6103), .sena
       (n_6088), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[3] [15]));
  CDN_flop \regs68H_reg[2][0] (.clk (\Clks[clk] ), .d (n_6111), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [0]));
  CDN_flop \regs68H_reg[2][1] (.clk (\Clks[clk] ), .d (n_6113), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [1]));
  CDN_flop \regs68H_reg[2][2] (.clk (\Clks[clk] ), .d (n_6114), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [2]));
  CDN_flop \regs68H_reg[2][3] (.clk (\Clks[clk] ), .d (n_6115), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [3]));
  CDN_flop \regs68H_reg[2][4] (.clk (\Clks[clk] ), .d (n_6116), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [4]));
  CDN_flop \regs68H_reg[2][5] (.clk (\Clks[clk] ), .d (n_6117), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [5]));
  CDN_flop \regs68H_reg[2][6] (.clk (\Clks[clk] ), .d (n_6118), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [6]));
  CDN_flop \regs68H_reg[2][7] (.clk (\Clks[clk] ), .d (n_6119), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [7]));
  CDN_flop \regs68H_reg[2][8] (.clk (\Clks[clk] ), .d (n_6120), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [8]));
  CDN_flop \regs68H_reg[2][9] (.clk (\Clks[clk] ), .d (n_6121), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [9]));
  CDN_flop \regs68H_reg[2][10] (.clk (\Clks[clk] ), .d (n_6122), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [10]));
  CDN_flop \regs68H_reg[2][11] (.clk (\Clks[clk] ), .d (n_6123), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [11]));
  CDN_flop \regs68H_reg[2][12] (.clk (\Clks[clk] ), .d (n_6124), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [12]));
  CDN_flop \regs68H_reg[2][13] (.clk (\Clks[clk] ), .d (n_6125), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [13]));
  CDN_flop \regs68H_reg[2][14] (.clk (\Clks[clk] ), .d (n_6126), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [14]));
  CDN_flop \regs68H_reg[2][15] (.clk (\Clks[clk] ), .d (n_6127), .sena
       (n_6112), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[2] [15]));
  CDN_flop \regs68H_reg[1][0] (.clk (\Clks[clk] ), .d (n_6135), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [0]));
  CDN_flop \regs68H_reg[1][1] (.clk (\Clks[clk] ), .d (n_6137), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [1]));
  CDN_flop \regs68H_reg[1][2] (.clk (\Clks[clk] ), .d (n_6138), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [2]));
  CDN_flop \regs68H_reg[1][3] (.clk (\Clks[clk] ), .d (n_6139), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [3]));
  CDN_flop \regs68H_reg[1][4] (.clk (\Clks[clk] ), .d (n_6140), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [4]));
  CDN_flop \regs68H_reg[1][5] (.clk (\Clks[clk] ), .d (n_6141), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [5]));
  CDN_flop \regs68H_reg[1][6] (.clk (\Clks[clk] ), .d (n_6142), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [6]));
  CDN_flop \regs68H_reg[1][7] (.clk (\Clks[clk] ), .d (n_6143), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [7]));
  CDN_flop \regs68H_reg[1][8] (.clk (\Clks[clk] ), .d (n_6144), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [8]));
  CDN_flop \regs68H_reg[1][9] (.clk (\Clks[clk] ), .d (n_6145), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [9]));
  CDN_flop \regs68H_reg[1][10] (.clk (\Clks[clk] ), .d (n_6146), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [10]));
  CDN_flop \regs68H_reg[1][11] (.clk (\Clks[clk] ), .d (n_6147), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [11]));
  CDN_flop \regs68H_reg[1][12] (.clk (\Clks[clk] ), .d (n_6148), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [12]));
  CDN_flop \regs68H_reg[1][13] (.clk (\Clks[clk] ), .d (n_6149), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [13]));
  CDN_flop \regs68H_reg[1][14] (.clk (\Clks[clk] ), .d (n_6150), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [14]));
  CDN_flop \regs68H_reg[1][15] (.clk (\Clks[clk] ), .d (n_6151), .sena
       (n_6136), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[1] [15]));
  CDN_flop \regs68H_reg[0][0] (.clk (\Clks[clk] ), .d (n_6159), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [0]));
  CDN_flop \regs68H_reg[0][1] (.clk (\Clks[clk] ), .d (n_6161), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [1]));
  CDN_flop \regs68H_reg[0][2] (.clk (\Clks[clk] ), .d (n_6162), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [2]));
  CDN_flop \regs68H_reg[0][3] (.clk (\Clks[clk] ), .d (n_6163), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [3]));
  CDN_flop \regs68H_reg[0][4] (.clk (\Clks[clk] ), .d (n_6164), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [4]));
  CDN_flop \regs68H_reg[0][5] (.clk (\Clks[clk] ), .d (n_6165), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [5]));
  CDN_flop \regs68H_reg[0][6] (.clk (\Clks[clk] ), .d (n_6166), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [6]));
  CDN_flop \regs68H_reg[0][7] (.clk (\Clks[clk] ), .d (n_6167), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [7]));
  CDN_flop \regs68H_reg[0][8] (.clk (\Clks[clk] ), .d (n_6168), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [8]));
  CDN_flop \regs68H_reg[0][9] (.clk (\Clks[clk] ), .d (n_6169), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [9]));
  CDN_flop \regs68H_reg[0][10] (.clk (\Clks[clk] ), .d (n_6170), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [10]));
  CDN_flop \regs68H_reg[0][11] (.clk (\Clks[clk] ), .d (n_6171), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [11]));
  CDN_flop \regs68H_reg[0][12] (.clk (\Clks[clk] ), .d (n_6172), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [12]));
  CDN_flop \regs68H_reg[0][13] (.clk (\Clks[clk] ), .d (n_6173), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [13]));
  CDN_flop \regs68H_reg[0][14] (.clk (\Clks[clk] ), .d (n_6174), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [14]));
  CDN_flop \regs68H_reg[0][15] (.clk (\Clks[clk] ), .d (n_6175), .sena
       (n_6160), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (\regs68H[0] [15]));
  CDN_flop \PcL_reg[0] (.clk (\Clks[clk] ), .d (n_6182), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[0]));
  CDN_flop \PcL_reg[1] (.clk (\Clks[clk] ), .d (n_6184), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[1]));
  CDN_flop \PcL_reg[2] (.clk (\Clks[clk] ), .d (n_6185), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[2]));
  CDN_flop \PcL_reg[3] (.clk (\Clks[clk] ), .d (n_6186), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[3]));
  CDN_flop \PcL_reg[4] (.clk (\Clks[clk] ), .d (n_6187), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[4]));
  CDN_flop \PcL_reg[5] (.clk (\Clks[clk] ), .d (n_6188), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[5]));
  CDN_flop \PcL_reg[6] (.clk (\Clks[clk] ), .d (n_6189), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[6]));
  CDN_flop \PcL_reg[7] (.clk (\Clks[clk] ), .d (n_6190), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[7]));
  CDN_flop \PcL_reg[8] (.clk (\Clks[clk] ), .d (n_6191), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[8]));
  CDN_flop \PcL_reg[9] (.clk (\Clks[clk] ), .d (n_6192), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[9]));
  CDN_flop \PcL_reg[10] (.clk (\Clks[clk] ), .d (n_6193), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[10]));
  CDN_flop \PcL_reg[11] (.clk (\Clks[clk] ), .d (n_6194), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[11]));
  CDN_flop \PcL_reg[12] (.clk (\Clks[clk] ), .d (n_6195), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[12]));
  CDN_flop \PcL_reg[13] (.clk (\Clks[clk] ), .d (n_6196), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[13]));
  CDN_flop \PcL_reg[14] (.clk (\Clks[clk] ), .d (n_6197), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[14]));
  CDN_flop \PcL_reg[15] (.clk (\Clks[clk] ), .d (n_6198), .sena
       (n_6183), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcL[15]));
  CDN_flop \PcH_reg[0] (.clk (\Clks[clk] ), .d (n_6205), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[0]));
  CDN_flop \PcH_reg[1] (.clk (\Clks[clk] ), .d (n_6207), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[1]));
  CDN_flop \PcH_reg[2] (.clk (\Clks[clk] ), .d (n_6208), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[2]));
  CDN_flop \PcH_reg[3] (.clk (\Clks[clk] ), .d (n_6209), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[3]));
  CDN_flop \PcH_reg[4] (.clk (\Clks[clk] ), .d (n_6210), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[4]));
  CDN_flop \PcH_reg[5] (.clk (\Clks[clk] ), .d (n_6211), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[5]));
  CDN_flop \PcH_reg[6] (.clk (\Clks[clk] ), .d (n_6212), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[6]));
  CDN_flop \PcH_reg[7] (.clk (\Clks[clk] ), .d (n_6213), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[7]));
  CDN_flop \PcH_reg[8] (.clk (\Clks[clk] ), .d (n_6214), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[8]));
  CDN_flop \PcH_reg[9] (.clk (\Clks[clk] ), .d (n_6215), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[9]));
  CDN_flop \PcH_reg[10] (.clk (\Clks[clk] ), .d (n_6216), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[10]));
  CDN_flop \PcH_reg[11] (.clk (\Clks[clk] ), .d (n_6217), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[11]));
  CDN_flop \PcH_reg[12] (.clk (\Clks[clk] ), .d (n_6218), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[12]));
  CDN_flop \PcH_reg[13] (.clk (\Clks[clk] ), .d (n_6219), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[13]));
  CDN_flop \PcH_reg[14] (.clk (\Clks[clk] ), .d (n_6220), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[14]));
  CDN_flop \PcH_reg[15] (.clk (\Clks[clk] ), .d (n_6221), .sena
       (n_6206), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (PcH[15]));
  CDN_flop \Ath_reg[0] (.clk (\Clks[clk] ), .d (n_6225), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[0]));
  CDN_flop \Ath_reg[1] (.clk (\Clks[clk] ), .d (n_6227), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[1]));
  CDN_flop \Ath_reg[2] (.clk (\Clks[clk] ), .d (n_6228), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[2]));
  CDN_flop \Ath_reg[3] (.clk (\Clks[clk] ), .d (n_6229), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[3]));
  CDN_flop \Ath_reg[4] (.clk (\Clks[clk] ), .d (n_6230), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[4]));
  CDN_flop \Ath_reg[5] (.clk (\Clks[clk] ), .d (n_6231), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[5]));
  CDN_flop \Ath_reg[6] (.clk (\Clks[clk] ), .d (n_6232), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[6]));
  CDN_flop \Ath_reg[7] (.clk (\Clks[clk] ), .d (n_6233), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[7]));
  CDN_flop \Ath_reg[8] (.clk (\Clks[clk] ), .d (n_6234), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[8]));
  CDN_flop \Ath_reg[9] (.clk (\Clks[clk] ), .d (n_6235), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[9]));
  CDN_flop \Ath_reg[10] (.clk (\Clks[clk] ), .d (n_6236), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[10]));
  CDN_flop \Ath_reg[11] (.clk (\Clks[clk] ), .d (n_6237), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[11]));
  CDN_flop \Ath_reg[12] (.clk (\Clks[clk] ), .d (n_6238), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[12]));
  CDN_flop \Ath_reg[13] (.clk (\Clks[clk] ), .d (n_6239), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[13]));
  CDN_flop \Ath_reg[14] (.clk (\Clks[clk] ), .d (n_6240), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[14]));
  CDN_flop \Ath_reg[15] (.clk (\Clks[clk] ), .d (n_6241), .sena
       (n_6226), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Ath[15]));
  CDN_flop \Atl_reg[0] (.clk (\Clks[clk] ), .d (n_6245), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[0]));
  CDN_flop \Atl_reg[1] (.clk (\Clks[clk] ), .d (n_6247), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[1]));
  CDN_flop \Atl_reg[2] (.clk (\Clks[clk] ), .d (n_6248), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[2]));
  CDN_flop \Atl_reg[3] (.clk (\Clks[clk] ), .d (n_6249), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[3]));
  CDN_flop \Atl_reg[4] (.clk (\Clks[clk] ), .d (n_6250), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[4]));
  CDN_flop \Atl_reg[5] (.clk (\Clks[clk] ), .d (n_6251), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[5]));
  CDN_flop \Atl_reg[6] (.clk (\Clks[clk] ), .d (n_6252), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[6]));
  CDN_flop \Atl_reg[7] (.clk (\Clks[clk] ), .d (n_6253), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[7]));
  CDN_flop \Atl_reg[8] (.clk (\Clks[clk] ), .d (n_6254), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[8]));
  CDN_flop \Atl_reg[9] (.clk (\Clks[clk] ), .d (n_6255), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[9]));
  CDN_flop \Atl_reg[10] (.clk (\Clks[clk] ), .d (n_6256), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[10]));
  CDN_flop \Atl_reg[11] (.clk (\Clks[clk] ), .d (n_6257), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[11]));
  CDN_flop \Atl_reg[12] (.clk (\Clks[clk] ), .d (n_6258), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[12]));
  CDN_flop \Atl_reg[13] (.clk (\Clks[clk] ), .d (n_6259), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[13]));
  CDN_flop \Atl_reg[14] (.clk (\Clks[clk] ), .d (n_6260), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[14]));
  CDN_flop \Atl_reg[15] (.clk (\Clks[clk] ), .d (n_6261), .sena
       (n_6246), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (Atl[15]));
  CDN_flop Pcl2Dbl_reg(.clk (\Clks[clk] ), .d (n_505), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (Pcl2Dbl));
  CDN_flop Pch2Dbh_reg(.clk (\Clks[clk] ), .d (n_644), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (Pch2Dbh));
  CDN_flop Pcl2Abl_reg(.clk (\Clks[clk] ), .d (n_537), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (Pcl2Abl));
  CDN_flop Pch2Abh_reg(.clk (\Clks[clk] ), .d (n_639), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (Pch2Abh));
  CDN_flop dbl2Pcl_reg(.clk (\Clks[clk] ), .d (n_554), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (dbl2Pcl));
  CDN_flop dbh2Pch_reg(.clk (\Clks[clk] ), .d (n_641), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (dbh2Pch));
  CDN_flop abh2Pch_reg(.clk (\Clks[clk] ), .d (n_1027), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (abh2Pch));
  CDN_flop abl2Pcl_reg(.clk (\Clks[clk] ), .d (n_555), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b0), .q (abl2Pcl));
  nor g2481 (n_8229, prenLatch[15], prenLatch[14], prenLatch[13],
       prenLatch[12]);
  nor g2482 (n_8230, prenLatch[11], prenLatch[10], prenLatch[9],
       prenLatch[8]);
  nor g2483 (n_8231, prenLatch[7], prenLatch[6], prenLatch[5],
       prenLatch[4]);
  nor g2484 (n_8232, prenLatch[3], prenLatch[2], prenLatch[1],
       prenLatch[0]);
  nand g2485 (n_8233, n_8229, n_8230, n_8231, n_8232);
  not g2486 (prenEmpty, n_8233);
  nor g2487 (n_439, n_8234, n_8235);
  nand g2488 (n_8234, prHbit[0], prHbit[3]);
  nand g2489 (n_8235, prHbit[1], prHbit[2]);
  nor g2490 (n_438, n_8235, n_8236);
  nor g2491 (n_437, n_8234, n_8237);
  nor g2492 (n_436, n_8236, n_8237);
  nor g2493 (n_435, n_8234, n_8238);
  nor g2494 (n_434, n_8236, n_8238);
  nor g2495 (n_433, n_8234, n_8239);
  nor g2496 (n_432, n_8236, n_8239);
  nor g2497 (n_431, n_8235, n_8240);
  nor g2498 (n_430, n_8235, n_8241);
  nor g2499 (n_429, n_8240, n_8237);
  nor g2500 (n_428, n_8241, n_8237);
  nor g2501 (n_427, n_8240, n_8238);
  nor g2502 (n_426, n_8241, n_8238);
  nor g2503 (n_424, n_8240, n_8239);
  nor g2504 (n_423, n_8241, n_8239);
  not g2505 (n_8242, prHbit[3]);
  not g2506 (n_8243, prHbit[0]);
  not g2507 (n_8244, prHbit[2]);
  not g2508 (n_8245, prHbit[1]);
  nand g2509 (n_8236, prHbit[3], n_8243);
  nand g2510 (n_8237, prHbit[2], n_8245);
  nand g2511 (n_8238, n_8244, prHbit[1]);
  nand g2512 (n_8239, n_8244, n_8245);
  nand g2513 (n_8240, n_8242, prHbit[0]);
  nand g2514 (n_8241, n_8242, n_8243);
  CDN_flop \movemRx_reg[0] (.clk (\Clks[clk] ), .d (n_6263), .sena
       (n_6264), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (movemRx[0]));
  CDN_flop \movemRx_reg[1] (.clk (\Clks[clk] ), .d (n_6265), .sena
       (n_6264), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (movemRx[1]));
  CDN_flop \movemRx_reg[2] (.clk (\Clks[clk] ), .d (n_6266), .sena
       (n_6264), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (movemRx[2]));
  CDN_flop \movemRx_reg[3] (.clk (\Clks[clk] ), .d (n_6267), .sena
       (n_6264), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (movemRx[3]));
  CDN_flop \prenLatch_reg[0] (.clk (\Clks[clk] ), .d (n_6269), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[0]));
  CDN_flop \prenLatch_reg[1] (.clk (\Clks[clk] ), .d (n_6271), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[1]));
  CDN_flop \prenLatch_reg[2] (.clk (\Clks[clk] ), .d (n_6272), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[2]));
  CDN_flop \prenLatch_reg[3] (.clk (\Clks[clk] ), .d (n_6273), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[3]));
  CDN_flop \prenLatch_reg[4] (.clk (\Clks[clk] ), .d (n_6274), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[4]));
  CDN_flop \prenLatch_reg[5] (.clk (\Clks[clk] ), .d (n_6275), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[5]));
  CDN_flop \prenLatch_reg[6] (.clk (\Clks[clk] ), .d (n_6276), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[6]));
  CDN_flop \prenLatch_reg[7] (.clk (\Clks[clk] ), .d (n_6277), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[7]));
  CDN_flop \prenLatch_reg[8] (.clk (\Clks[clk] ), .d (n_6278), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[8]));
  CDN_flop \prenLatch_reg[9] (.clk (\Clks[clk] ), .d (n_6279), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[9]));
  CDN_flop \prenLatch_reg[10] (.clk (\Clks[clk] ), .d (n_6280), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[10]));
  CDN_flop \prenLatch_reg[11] (.clk (\Clks[clk] ), .d (n_6281), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[11]));
  CDN_flop \prenLatch_reg[12] (.clk (\Clks[clk] ), .d (n_6282), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[12]));
  CDN_flop \prenLatch_reg[13] (.clk (\Clks[clk] ), .d (n_6283), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[13]));
  CDN_flop \prenLatch_reg[14] (.clk (\Clks[clk] ), .d (n_6284), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[14]));
  CDN_flop \prenLatch_reg[15] (.clk (\Clks[clk] ), .d (n_6285), .sena
       (n_6270), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (prenLatch[15]));
  CDN_flop dcr4_reg(.clk (\Clks[clk] ), .d (Abd[4]), .sena (n_643),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd (1'b0),
       .q (dcr4));
  CDN_flop \dcrOutput_reg[0] (.clk (\Clks[clk] ), .d (dcrCode[0]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[0]));
  CDN_flop \dcrOutput_reg[1] (.clk (\Clks[clk] ), .d (dcrCode[1]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[1]));
  CDN_flop \dcrOutput_reg[2] (.clk (\Clks[clk] ), .d (dcrCode[2]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[2]));
  CDN_flop \dcrOutput_reg[3] (.clk (\Clks[clk] ), .d (dcrCode[3]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[3]));
  CDN_flop \dcrOutput_reg[4] (.clk (\Clks[clk] ), .d (dcrCode[4]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[4]));
  CDN_flop \dcrOutput_reg[5] (.clk (\Clks[clk] ), .d (dcrCode[5]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[5]));
  CDN_flop \dcrOutput_reg[6] (.clk (\Clks[clk] ), .d (dcrCode[6]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[6]));
  CDN_flop \dcrOutput_reg[7] (.clk (\Clks[clk] ), .d (dcrCode[7]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[7]));
  CDN_flop \dcrOutput_reg[8] (.clk (\Clks[clk] ), .d (dcrCode[8]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[8]));
  CDN_flop \dcrOutput_reg[9] (.clk (\Clks[clk] ), .d (dcrCode[9]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[9]));
  CDN_flop \dcrOutput_reg[10] (.clk (\Clks[clk] ), .d (dcrCode[10]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[10]));
  CDN_flop \dcrOutput_reg[11] (.clk (\Clks[clk] ), .d (dcrCode[11]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[11]));
  CDN_flop \dcrOutput_reg[12] (.clk (\Clks[clk] ), .d (dcrCode[12]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[12]));
  CDN_flop \dcrOutput_reg[13] (.clk (\Clks[clk] ), .d (dcrCode[13]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[13]));
  CDN_flop \dcrOutput_reg[14] (.clk (\Clks[clk] ), .d (dcrCode[14]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[14]));
  CDN_flop \dcrOutput_reg[15] (.clk (\Clks[clk] ), .d (dcrCode[15]),
       .sena (n_6287), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (dcrOutput[15]));
  CDN_flop \alub_reg[0] (.clk (\Clks[clk] ), .d (n_6291), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[0]));
  CDN_flop \alub_reg[1] (.clk (\Clks[clk] ), .d (n_6293), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[1]));
  CDN_flop \alub_reg[2] (.clk (\Clks[clk] ), .d (n_6294), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[2]));
  CDN_flop \alub_reg[3] (.clk (\Clks[clk] ), .d (n_6295), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[3]));
  CDN_flop \alub_reg[4] (.clk (\Clks[clk] ), .d (n_6296), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[4]));
  CDN_flop \alub_reg[5] (.clk (\Clks[clk] ), .d (n_6297), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[5]));
  CDN_flop \alub_reg[6] (.clk (\Clks[clk] ), .d (n_6298), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[6]));
  CDN_flop \alub_reg[7] (.clk (\Clks[clk] ), .d (n_6299), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[7]));
  CDN_flop \alub_reg[8] (.clk (\Clks[clk] ), .d (n_6300), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[8]));
  CDN_flop \alub_reg[9] (.clk (\Clks[clk] ), .d (n_6301), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[9]));
  CDN_flop \alub_reg[10] (.clk (\Clks[clk] ), .d (n_6302), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[10]));
  CDN_flop \alub_reg[11] (.clk (\Clks[clk] ), .d (n_6303), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[11]));
  CDN_flop \alub_reg[12] (.clk (\Clks[clk] ), .d (n_6304), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[12]));
  CDN_flop \alub_reg[13] (.clk (\Clks[clk] ), .d (n_6305), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[13]));
  CDN_flop \alub_reg[14] (.clk (\Clks[clk] ), .d (n_6306), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[14]));
  CDN_flop \alub_reg[15] (.clk (\Clks[clk] ), .d (n_6307), .sena
       (n_6292), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0),
       .q (alub[15]));
  nor g2569 (dobIdle, \Nanod[dobCtrl] [0], \Nanod[dobCtrl] [1]);
  and g2570 (n_10, n_9, pswS);
  not g2571 (n_6349, pswS);
  and g2572 (n_11, n_6349, n_9);
  or g2574 (n_16, \Irdecod[rxIsUsp] , \Nanod[ssp] );
  or g2 (n_19, n_8, n_16);
  not g2575 (n_17, \Nanod[ssp] );
  and g2576 (n_492, n_17, \Irdecod[rxIsUsp] );
  not g5 (n_18, n_16);
  and g2577 (n_493, n_18, n_8);
  not g2578 (n_20, n_19);
  and g2579 (n_494, n_20, n_9);
  nor g2584 (n_495, \Nanod[ssp] , \Irdecod[rxIsUsp] , n_8, n_9);
  and g2594 (n_501, n_20, n_10);
  nor g18 (n_32, \Nanod[ssp] , \Irdecod[rxIsUsp] , n_8, n_10);
  not g19 (n_33, n_11);
  nand g2598 (n_34, n_32, n_33);
  not g2599 (n_503, n_34);
  nor g2606 (n_29, rxl2Dbl, ryl2Dbl, \Nanod[ftu2Dbl] , \Nanod[au2Db] );
  nor g2607 (n_28, \Nanod[atl2Dbl] , Pcl2Dbl);
  nand g2608 (n_30, n_28, n_29);
  not g2609 (n_517, n_30);
  nor g2614 (n_535, ryl2Abd, rxl2Abd, \Nanod[dbin2Abd] ,
       \Nanod[alu2Abd] );
  nor g2622 (n_8375, Pcl2Abl, rxl2Abl, ryl2Abl, \Nanod[ftu2Abl] );
  nor g2623 (n_8374, \Nanod[au2Ab] , \Nanod[aob2Ab] , \Nanod[atl2Abl] );
  nand g2624 (n_8376, n_8374, n_8375);
  not g2625 (n_551, n_8376);
  nor g2631 (n_8377, \Nanod[rxh2dbh] , \Nanod[ryh2dbh] , \Nanod[au2Db]
       , \Nanod[ath2Dbh] );
  not g2632 (n_8378, Pch2Dbh);
  nand g2633 (n_8379, n_8377, n_8378);
  not g2634 (n_653, n_8379);
  nor g2641 (n_8381, Pch2Abh, \Nanod[rxh2abh] , \Nanod[ryh2abh] ,
       \Nanod[au2Ab] );
  nor g2642 (n_8380, \Nanod[aob2Ab] , \Nanod[ath2Abh] );
  nand g2643 (n_8382, n_8380, n_8381);
  not g2644 (n_666, n_8382);
  nor g2645 (n_669, n_207, n_8386);
  nand g2646 (n_207, n_205, n_206);
  not g2647 (n_205, actualRy[0]);
  not g2648 (n_206, actualRy[3]);
  nand g2649 (n_8386, n_8384, n_8385);
  not g2650 (n_8384, actualRy[1]);
  nor g2651 (n_8385, actualRy[4], actualRy[2]);
  nor g2652 (n_719, n_8386, n_13);
  nand g2653 (n_13, actualRy[0], n_206);
  nor g2654 (n_737, n_207, n_15);
  nand g2655 (n_15, n_8385, actualRy[1]);
  nor g2656 (n_755, n_15, n_13);
  nor g2657 (n_773, n_207, n_8389);
  nand g2658 (n_8389, n_8384, n_8388);
  nor g2659 (n_8388, actualRy[4], n_8387);
  not g2660 (n_8387, actualRy[2]);
  nor g2661 (n_791, n_8389, n_13);
  nor g2662 (n_809, n_207, n_8390);
  nand g2663 (n_8390, n_8388, actualRy[1]);
  nor g2664 (n_827, n_8390, n_13);
  nor g2665 (n_845, n_8386, n_8391);
  nand g2666 (n_8391, n_205, actualRy[3]);
  nor g2667 (n_863, n_8386, n_8392);
  nand g2668 (n_8392, actualRy[0], actualRy[3]);
  nor g2669 (n_881, n_15, n_8391);
  nor g2670 (n_899, n_15, n_8392);
  nor g2671 (n_917, n_8389, n_8391);
  nor g2672 (n_935, n_8389, n_8392);
  nor g2673 (n_953, n_8390, n_8391);
  nor g2674 (n_971, n_8390, n_8392);
  nor g2675 (n_989, n_207, n_38);
  nand g2676 (n_38, n_8384, n_37);
  nor g2677 (n_37, n_36, actualRy[2]);
  not g2678 (n_36, actualRy[4]);
  nor g2679 (n_1007, n_38, n_13);
  nor g2775 (n_8444, ryl2Dbd, rxl2Dbd, \Nanod[alue2Dbd] ,
       \Nanod[dbin2Dbd] );
  nor g2776 (n_8443, \Nanod[alu2Dbd] , \Nanod[dcr2Dbd] );
  nand g2777 (n_8445, n_8443, n_8444);
  not g2778 (n_1357, n_8445);
  nand g2870 (n_6, n_8502, n_8503, n_8504, n_208);
  nor g2871 (n_5664, n_6, actualRx[0]);
  nor g2872 (n_5585, n_6, n_209);
  nand g2873 (n_8505, n_8502, n_8503, n_8504, actualRx[1]);
  nor g2874 (n_5506, n_8505, actualRx[0]);
  nor g2875 (n_5427, n_8505, n_209);
  nand g2876 (n_8506, n_8502, n_8503, actualRx[2], n_208);
  nor g2877 (n_5348, n_8506, actualRx[0]);
  nor g2878 (n_5269, n_8506, n_209);
  nand g2879 (n_8507, n_8502, n_8503, actualRx[2], actualRx[1]);
  nor g2880 (n_5190, n_8507, actualRx[0]);
  nor g2881 (n_5111, n_8507, n_209);
  nand g2882 (n_62, n_8502, actualRx[3], n_8504, n_208);
  nor g2883 (n_5032, n_62, actualRx[0]);
  nor g2884 (n_4953, n_62, n_209);
  nand g2885 (n_76, n_8502, actualRx[3], n_8504, actualRx[1]);
  nor g2886 (n_4874, n_76, actualRx[0]);
  nor g2887 (n_4795, n_76, n_209);
  nand g2888 (n_90, n_8502, actualRx[3], actualRx[2], n_208);
  nor g2889 (n_4716, n_90, actualRx[0]);
  nor g42 (n_4637, n_90, n_209);
  nand g43 (n_210, n_8502, actualRx[3], actualRx[2], actualRx[1]);
  nor g45 (n_4558, n_210, actualRx[0]);
  nor g48 (n_4479, n_210, n_209);
  nand g49 (n_118, actualRx[4], n_8503, n_8504, n_208);
  nor g51 (n_4400, n_118, actualRx[0]);
  not g53 (n_209, actualRx[0]);
  nor g2890 (n_4315, n_118, n_209);
  not g63 (n_8502, actualRx[4]);
  not g2895 (n_8503, actualRx[3]);
  not g2896 (n_8504, actualRx[2]);
  not g2897 (n_208, actualRx[1]);
  and g3078 (n_502, n_8616, n_8617, n_8618, n_11);
  not g3079 (n_8616, n_10);
  not g3080 (n_8617, n_8);
  not g3081 (n_8618, n_16);
endmodule

module fx68k_or_op_1324(A, Z);
  input [1:0] A;
  output Z;
  wire [1:0] A;
  wire Z;
  wire n_3;
  nor g1 (n_3, A[0], A[1]);
  not g2 (Z, n_3);
endmodule

module fx68k_or_op_1325(A, Z);
  input [1:0] A;
  output Z;
  wire [1:0] A;
  wire Z;
  wire n_3;
  nor g1 (n_3, A[0], A[1]);
  not g2 (Z, n_3);
endmodule

module fx68k_nDecoder3(\Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] ,
     \Clks[extReset] , \Clks[clk] , \Irdecod[inhibitCcr] ,
     \Irdecod[macroTvn] , \Irdecod[ftuConst] , \Irdecod[ryIsAreg] ,
     \Irdecod[rxIsAreg] , \Irdecod[ry] , \Irdecod[rx] ,
     \Irdecod[isMovep] , \Irdecod[isByte] , \Irdecod[movemPreDecr] ,
     \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] ,
     \Irdecod[rxIsDt] , \Irdecod[toCcr] , \Irdecod[implicitSp] ,
     \Irdecod[isTas] , \Irdecod[isPcRel] , \Nanod[abdIsByte] ,
     \Nanod[dblDbh] , \Nanod[dblDbd] , \Nanod[ablAbh] , \Nanod[ablAbd]
     , \Nanod[extAbh] , \Nanod[extDbh] , \Nanod[dbin2Dbd] ,
     \Nanod[dbin2Abd] , \Nanod[au2Pc] , \Nanod[au2Ab] , \Nanod[au2Db] ,
     \Nanod[alu2Abd] , \Nanod[alu2Dbd] , \Nanod[abd2Alub] ,
     \Nanod[dbd2Alub] , \Nanod[alue2Dbd] , \Nanod[dbd2Alue] ,
     \Nanod[dcr2Dbd] , \Nanod[abd2Dcr] , \Nanod[aluFinish] ,
     \Nanod[aluInit] , \Nanod[aluActrl] , \Nanod[aluDctrl] ,
     \Nanod[aluColumn] , \Nanod[rxlDbl] , \Nanod[rz] , \Nanod[abl2ryl]
     , \Nanod[dbl2ryl] , \Nanod[ryh2abh] , \Nanod[ryh2dbh] ,
     \Nanod[ryl2ab] , \Nanod[ryl2db] , \Nanod[abh2ryh] ,
     \Nanod[dbh2ryh] , \Nanod[abh2rxh] , \Nanod[abl2rxl] ,
     \Nanod[rxl2ab] , \Nanod[rxl2db] , \Nanod[dbh2rxh] ,
     \Nanod[dbl2rxl] , \Nanod[rxh2abh] , \Nanod[rxh2dbh] ,
     \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl] , \Nanod[pchdbh]
     , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl] ,
     \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
     \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
     \Nanod[dobCtrl] , \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob]
     , \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
     \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
     \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
     \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] , \Nanod[auCntrl]
     , \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
     \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
     \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
     \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
     \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
     \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
     \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
     \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
     \Nanod[waitBusFinish] , \Nanod[permStart] , enT2, enT4,
     microLatch, nanoLatch);
  input \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset]
       , \Clks[clk] , \Irdecod[inhibitCcr] , \Irdecod[ryIsAreg] ,
       \Irdecod[rxIsAreg] , \Irdecod[isMovep] , \Irdecod[isByte] ,
       \Irdecod[movemPreDecr] , \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp]
       , \Irdecod[ryIsDt] , \Irdecod[rxIsDt] , \Irdecod[toCcr] ,
       \Irdecod[implicitSp] , \Irdecod[isTas] , \Irdecod[isPcRel] ,
       enT2, enT4;
  input [5:0] \Irdecod[macroTvn] ;
  input [15:0] \Irdecod[ftuConst] ;
  input [2:0] \Irdecod[ry] , \Irdecod[rx] ;
  input [16:0] microLatch;
  input [67:0] nanoLatch;
  output \Nanod[abdIsByte] , \Nanod[dblDbh] , \Nanod[dblDbd] ,
       \Nanod[ablAbh] , \Nanod[ablAbd] , \Nanod[extAbh] ,
       \Nanod[extDbh] , \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] ,
       \Nanod[au2Pc] , \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd]
       , \Nanod[alu2Dbd] , \Nanod[abd2Alub] , \Nanod[dbd2Alub] ,
       \Nanod[alue2Dbd] , \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] ,
       \Nanod[abd2Dcr] , \Nanod[aluFinish] , \Nanod[aluInit] ,
       \Nanod[aluActrl] , \Nanod[rxlDbl] , \Nanod[rz] , \Nanod[abl2ryl]
       , \Nanod[dbl2ryl] , \Nanod[ryh2abh] , \Nanod[ryh2dbh] ,
       \Nanod[ryl2ab] , \Nanod[ryl2db] , \Nanod[abh2ryh] ,
       \Nanod[dbh2ryh] , \Nanod[abh2rxh] , \Nanod[abl2rxl] ,
       \Nanod[rxl2ab] , \Nanod[rxl2db] , \Nanod[dbh2rxh] ,
       \Nanod[dbl2rxl] , \Nanod[rxh2abh] , \Nanod[rxh2dbh] ,
       \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl] ,
       \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
       , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
       \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
       \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob] ,
       \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
       \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
       \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
       \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] ,
       \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
       \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
       \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
       \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
       \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
       \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
       \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
       \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
       \Nanod[waitBusFinish] , \Nanod[permStart] ;
  output [1:0] \Nanod[aluDctrl] , \Nanod[dobCtrl] ;
  output [2:0] \Nanod[aluColumn] , \Nanod[auCntrl] ;
  wire \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset] ,
       \Clks[clk] , \Irdecod[inhibitCcr] , \Irdecod[ryIsAreg] ,
       \Irdecod[rxIsAreg] , \Irdecod[isMovep] , \Irdecod[isByte] ,
       \Irdecod[movemPreDecr] , \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp]
       , \Irdecod[ryIsDt] , \Irdecod[rxIsDt] , \Irdecod[toCcr] ,
       \Irdecod[implicitSp] , \Irdecod[isTas] , \Irdecod[isPcRel] ,
       enT2, enT4;
  wire [5:0] \Irdecod[macroTvn] ;
  wire [15:0] \Irdecod[ftuConst] ;
  wire [2:0] \Irdecod[ry] , \Irdecod[rx] ;
  wire [16:0] microLatch;
  wire [67:0] nanoLatch;
  wire \Nanod[abdIsByte] , \Nanod[dblDbh] , \Nanod[dblDbd] ,
       \Nanod[ablAbh] , \Nanod[ablAbd] , \Nanod[extAbh] ,
       \Nanod[extDbh] , \Nanod[dbin2Dbd] , \Nanod[dbin2Abd] ,
       \Nanod[au2Pc] , \Nanod[au2Ab] , \Nanod[au2Db] , \Nanod[alu2Abd]
       , \Nanod[alu2Dbd] , \Nanod[abd2Alub] , \Nanod[dbd2Alub] ,
       \Nanod[alue2Dbd] , \Nanod[dbd2Alue] , \Nanod[dcr2Dbd] ,
       \Nanod[abd2Dcr] , \Nanod[aluFinish] , \Nanod[aluInit] ,
       \Nanod[aluActrl] , \Nanod[rxlDbl] , \Nanod[rz] , \Nanod[abl2ryl]
       , \Nanod[dbl2ryl] , \Nanod[ryh2abh] , \Nanod[ryh2dbh] ,
       \Nanod[ryl2ab] , \Nanod[ryl2db] , \Nanod[abh2ryh] ,
       \Nanod[dbh2ryh] , \Nanod[abh2rxh] , \Nanod[abl2rxl] ,
       \Nanod[rxl2ab] , \Nanod[rxl2db] , \Nanod[dbh2rxh] ,
       \Nanod[dbl2rxl] , \Nanod[rxh2abh] , \Nanod[rxh2dbh] ,
       \Nanod[pchabh] , \Nanod[pclabl] , \Nanod[pcldbl] ,
       \Nanod[pchdbh] , \Nanod[ssp] , \Nanod[reg2dbh] , \Nanod[reg2dbl]
       , \Nanod[dbl2reg] , \Nanod[dbh2reg] , \Nanod[reg2abh] ,
       \Nanod[reg2abl] , \Nanod[abl2reg] , \Nanod[abh2reg] ,
       \Nanod[updSsw] , \Nanod[aob2Ab] , \Nanod[au2Aob] ,
       \Nanod[ab2Aob] , \Nanod[db2Aob] , \Nanod[ath2Abh] ,
       \Nanod[ath2Dbh] , \Nanod[dbh2Ath] , \Nanod[abh2Ath] ,
       \Nanod[atl2Dbl] , \Nanod[atl2Abl] , \Nanod[abl2Atl] ,
       \Nanod[dbl2Atl] , \Nanod[toIrc] , \Nanod[todbin] ,
       \Nanod[noSpAlign] , \Nanod[auClkEn] , \Nanod[Ir2Ird] ,
       \Nanod[initST] , \Nanod[ssw2Ftu] , \Nanod[ird2Ftu] ,
       \Nanod[pswIToFtu] , \Nanod[ftu2Ccr] , \Nanod[sr2Ftu] ,
       \Nanod[ftu2Sr] , \Nanod[inl2psw] , \Nanod[updPren] ,
       \Nanod[abl2Pren] , \Nanod[ftu2Abl] , \Nanod[ftu2Dbl] ,
       \Nanod[const2Ftu] , \Nanod[tvn2Ftu] , \Nanod[clrTpend] ,
       \Nanod[updTpend] , \Nanod[noHighByte] , \Nanod[noLowByte] ,
       \Nanod[isRmc] , \Nanod[busByte] , \Nanod[isWrite] ,
       \Nanod[waitBusFinish] , \Nanod[permStart] ;
  wire [1:0] \Nanod[aluDctrl] , \Nanod[dobCtrl] ;
  wire [2:0] \Nanod[aluColumn] , \Nanod[auCntrl] ;
  wire [3:0] ftuCtrl;
  wire isPcRel, n_103, n_104, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_133;
  wire n_134, n_139, n_142, n_143, n_144, n_152, n_154, n_156;
  wire n_158, n_160, n_162, n_163, n_165, n_166, n_168, n_170;
  wire n_172, n_173, n_175, n_176, n_178, n_180, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_406;
  wire n_407, n_410, n_413, n_416, n_418, n_420, n_421, n_424;
  wire n_425, n_428, n_432, n_433, n_435, n_436, n_439, n_441;
  wire n_443, n_444, n_447, n_451, n_454, n_456, n_457, n_459;
  wire n_460, n_463, n_465, n_466, n_468, n_469, n_471, n_472;
  wire n_474, n_475, n_478, n_480, n_481, n_483, n_484, n_485;
  wire n_486, n_489, n_494, n_499, n_502, n_504, n_506, n_509;
  wire n_514, n_517, n_522, n_525, n_526, n_531, n_536, n_541;
  wire n_546, n_547, n_549, n_554, pcRelAbh, pcRelAbl, pcRelDbh,
       pcRelDbl;
  assign \Nanod[busByte]  = nanoLatch[42];
  assign \Nanod[noLowByte]  = nanoLatch[55];
  assign \Nanod[noHighByte]  = nanoLatch[54];
  assign \Nanod[updTpend]  = \Nanod[const2Ftu] ;
  assign \Nanod[Ir2Ird]  = nanoLatch[67];
  assign \Nanod[aob2Ab]  = \Nanod[updSsw] ;
  assign \Nanod[abh2reg]  = nanoLatch[7];
  assign \Nanod[abl2reg]  = nanoLatch[36];
  assign \Nanod[reg2abl]  = nanoLatch[37];
  assign \Nanod[reg2abh]  = nanoLatch[8];
  assign \Nanod[dbh2reg]  = nanoLatch[5];
  assign \Nanod[dbl2reg]  = nanoLatch[33];
  assign \Nanod[reg2dbl]  = nanoLatch[32];
  assign \Nanod[reg2dbh]  = nanoLatch[6];
  assign \Nanod[ssp]  = nanoLatch[24];
  assign \Nanod[rz]  = nanoLatch[43];
  assign \Nanod[rxlDbl]  = nanoLatch[40];
  assign \Nanod[aluColumn] [0] = nanoLatch[65];
  assign \Nanod[aluColumn] [1] = nanoLatch[64];
  assign \Nanod[aluColumn] [2] = nanoLatch[63];
  assign \Nanod[aluDctrl] [0] = nanoLatch[51];
  assign \Nanod[aluDctrl] [1] = nanoLatch[52];
  assign \Nanod[aluActrl]  = nanoLatch[50];
  assign \Nanod[dbin2Abd]  = nanoLatch[46];
  assign \Nanod[dbin2Dbd]  = nanoLatch[47];
  assign \Nanod[abdIsByte]  = nanoLatch[38];
  fx68k_or_op_1324 g36(.A (nanoLatch[4:3]), .Z (\Nanod[permStart] ));
  fx68k_or_op_1325 g37(.A ({nanoLatch[56], nanoLatch[53]}), .Z
       (\Nanod[isWrite] ));
  or g2 (n_123, n_103, n_104);
  or g33 (\Nanod[ftu2Dbl] , n_139, \Nanod[inl2psw] );
  or g34 (n_142, \Nanod[inl2psw] , \Nanod[clrTpend] );
  or g35 (\Nanod[initST] , n_142, n_143);
  or g38 (n_144, nanoLatch[66], nanoLatch[60]);
  or g39 (\Nanod[waitBusFinish] , n_144, \Nanod[isWrite] );
  and g45 (isPcRel, \Irdecod[isPcRel] , n_152);
  and g47 (pcRelDbl, isPcRel, n_154);
  and g49 (pcRelDbh, isPcRel, n_156);
  and g50 (pcRelAbl, isPcRel, nanoLatch[40]);
  and g51 (pcRelAbh, isPcRel, nanoLatch[22]);
  or g52 (\Nanod[pcldbl] , nanoLatch[39], pcRelDbl);
  or g53 (\Nanod[pchdbh] , n_158, pcRelDbh);
  or g54 (\Nanod[pclabl] , nanoLatch[41], pcRelAbl);
  or g55 (\Nanod[pchabh] , n_160, pcRelAbh);
  and g57 (n_163, nanoLatch[32], n_162);
  and g58 (n_202, n_163, nanoLatch[40]);
  and g60 (n_166, nanoLatch[37], n_165);
  and g61 (n_201, n_166, n_154);
  and g62 (n_168, nanoLatch[33], n_162);
  and g63 (n_204, n_168, nanoLatch[40]);
  and g64 (n_170, nanoLatch[36], n_165);
  and g65 (n_200, n_170, n_154);
  and g67 (n_173, nanoLatch[6], n_172);
  and g68 (n_206, n_173, nanoLatch[22]);
  and g70 (n_176, nanoLatch[8], n_175);
  and g71 (n_205, n_176, n_156);
  and g72 (n_178, nanoLatch[5], n_172);
  and g73 (n_203, n_178, nanoLatch[22]);
  and g74 (n_180, nanoLatch[7], n_175);
  and g75 (n_199, n_180, n_156);
  and g77 (n_198, n_178, n_156);
  and g79 (n_197, n_180, nanoLatch[22]);
  and g81 (n_192, n_168, n_154);
  and g83 (n_191, n_170, nanoLatch[40]);
  and g85 (n_196, n_163, n_154);
  and g87 (n_195, n_166, nanoLatch[40]);
  and g89 (n_194, n_173, n_156);
  and g91 (n_193, n_176, nanoLatch[22]);
  and g92 (n_207, \Irdecod[isTas] , nanoLatch[42]);
  not g1 (n_134, nanoLatch[19]);
  CDN_flop \Nanod_reg[dblDbh] (.clk (\Clks[clk] ), .d (nanoLatch[15]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[dblDbh] ));
  CDN_flop \Nanod_reg[dblDbd] (.clk (\Clks[clk] ), .d (nanoLatch[34]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[dblDbd] ));
  CDN_flop \Nanod_reg[ablAbh] (.clk (\Clks[clk] ), .d (nanoLatch[14]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[ablAbh] ));
  CDN_flop \Nanod_reg[ablAbd] (.clk (\Clks[clk] ), .d (nanoLatch[35]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[ablAbd] ));
  CDN_flop \Nanod_reg[extAbh] (.clk (\Clks[clk] ), .d (nanoLatch[13]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[extAbh] ));
  CDN_flop \Nanod_reg[extDbh] (.clk (\Clks[clk] ), .d (nanoLatch[12]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[extDbh] ));
  CDN_flop \Nanod_reg[alu2Abd] (.clk (\Clks[clk] ), .d (nanoLatch[45]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[alu2Abd] ));
  CDN_flop \Nanod_reg[alu2Dbd] (.clk (\Clks[clk] ), .d (nanoLatch[44]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[alu2Dbd] ));
  CDN_flop \Nanod_reg[abd2Alub] (.clk (\Clks[clk] ), .d
       (nanoLatch[48]), .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl
       (1'b0), .srd (1'b0), .q (\Nanod[abd2Alub] ));
  CDN_flop \Nanod_reg[dbd2Alub] (.clk (\Clks[clk] ), .d
       (nanoLatch[49]), .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl
       (1'b0), .srd (1'b0), .q (\Nanod[dbd2Alub] ));
  CDN_flop \Nanod_reg[alue2Dbd] (.clk (\Clks[clk] ), .d (n_116), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[alue2Dbd] ));
  CDN_flop \Nanod_reg[dbd2Alue] (.clk (\Clks[clk] ), .d (n_117), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dbd2Alue] ));
  CDN_flop \Nanod_reg[dcr2Dbd] (.clk (\Clks[clk] ), .d (n_118), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dcr2Dbd] ));
  CDN_flop \Nanod_reg[abd2Dcr] (.clk (\Clks[clk] ), .d (n_119), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[abd2Dcr] ));
  CDN_flop \Nanod_reg[dobCtrl][0] (.clk (\Clks[clk] ), .d
       (nanoLatch[53]), .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl
       (1'b0), .srd (1'b0), .q (\Nanod[dobCtrl] [0]));
  CDN_flop \Nanod_reg[dobCtrl][1] (.clk (\Clks[clk] ), .d
       (nanoLatch[56]), .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl
       (1'b0), .srd (1'b0), .q (\Nanod[dobCtrl] [1]));
  CDN_flop \Nanod_reg[aob2Ab] (.clk (\Clks[clk] ), .d (n_104), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[updSsw] ));
  CDN_flop \Nanod_reg[ath2Abh] (.clk (\Clks[clk] ), .d (n_120), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[ath2Abh] ));
  CDN_flop \Nanod_reg[ath2Dbh] (.clk (\Clks[clk] ), .d (n_121), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[ath2Dbh] ));
  CDN_flop \Nanod_reg[dbh2Ath] (.clk (\Clks[clk] ), .d (n_122), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dbh2Ath] ));
  CDN_flop \Nanod_reg[abh2Ath] (.clk (\Clks[clk] ), .d (n_123), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[abh2Ath] ));
  CDN_flop \Nanod_reg[atl2Dbl] (.clk (\Clks[clk] ), .d (n_124), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[atl2Dbl] ));
  CDN_flop \Nanod_reg[atl2Abl] (.clk (\Clks[clk] ), .d (n_125), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[atl2Abl] ));
  CDN_flop \Nanod_reg[abl2Atl] (.clk (\Clks[clk] ), .d (n_126), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[abl2Atl] ));
  CDN_flop \Nanod_reg[dbl2Atl] (.clk (\Clks[clk] ), .d (n_127), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dbl2Atl] ));
  CDN_flop \Nanod_reg[toIrc] (.clk (\Clks[clk] ), .d (nanoLatch[66]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[toIrc] ));
  CDN_flop \Nanod_reg[todbin] (.clk (\Clks[clk] ), .d (nanoLatch[60]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (\Nanod[todbin] ));
  CDN_flop \Nanod_reg[auCntrl][0] (.clk (\Clks[clk] ), .d
       (nanoLatch[16]), .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl
       (1'b0), .srd (1'b0), .q (\Nanod[auCntrl] [0]));
  CDN_flop \Nanod_reg[auCntrl][1] (.clk (\Clks[clk] ), .d
       (nanoLatch[17]), .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl
       (1'b0), .srd (1'b0), .q (\Nanod[auCntrl] [1]));
  CDN_flop \Nanod_reg[auCntrl][2] (.clk (\Clks[clk] ), .d
       (nanoLatch[18]), .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl
       (1'b0), .srd (1'b0), .q (\Nanod[auCntrl] [2]));
  CDN_flop \Nanod_reg[noSpAlign] (.clk (\Clks[clk] ), .d (n_133), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[noSpAlign] ));
  CDN_flop \Nanod_reg[auClkEn] (.clk (\Clks[clk] ), .d (n_134), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[auClkEn] ));
  CDN_flop \ftuCtrl_reg[0] (.clk (\Clks[clk] ), .d (nanoLatch[28]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (ftuCtrl[0]));
  CDN_flop \ftuCtrl_reg[1] (.clk (\Clks[clk] ), .d (nanoLatch[27]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (ftuCtrl[1]));
  CDN_flop \ftuCtrl_reg[2] (.clk (\Clks[clk] ), .d (nanoLatch[26]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (ftuCtrl[2]));
  CDN_flop \ftuCtrl_reg[3] (.clk (\Clks[clk] ), .d (nanoLatch[25]),
       .sena (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (ftuCtrl[3]));
  not g145 (n_152, nanoLatch[43]);
  not g146 (n_154, nanoLatch[40]);
  not g147 (n_156, nanoLatch[22]);
  not g148 (n_162, \Nanod[pcldbl] );
  not g149 (n_165, \Nanod[pclabl] );
  not g150 (n_172, \Nanod[pchdbh] );
  not g151 (n_175, \Nanod[pchabh] );
  CDN_flop \Nanod_reg[abl2ryl] (.clk (\Clks[clk] ), .d (n_191), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[abl2ryl] ));
  CDN_flop \Nanod_reg[dbl2ryl] (.clk (\Clks[clk] ), .d (n_192), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dbl2ryl] ));
  CDN_flop \Nanod_reg[ryh2abh] (.clk (\Clks[clk] ), .d (n_193), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[ryh2abh] ));
  CDN_flop \Nanod_reg[ryh2dbh] (.clk (\Clks[clk] ), .d (n_194), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[ryh2dbh] ));
  CDN_flop \Nanod_reg[ryl2ab] (.clk (\Clks[clk] ), .d (n_195), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[ryl2ab] ));
  CDN_flop \Nanod_reg[ryl2db] (.clk (\Clks[clk] ), .d (n_196), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[ryl2db] ));
  CDN_flop \Nanod_reg[abh2ryh] (.clk (\Clks[clk] ), .d (n_197), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[abh2ryh] ));
  CDN_flop \Nanod_reg[dbh2ryh] (.clk (\Clks[clk] ), .d (n_198), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dbh2ryh] ));
  CDN_flop \Nanod_reg[abh2rxh] (.clk (\Clks[clk] ), .d (n_199), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[abh2rxh] ));
  CDN_flop \Nanod_reg[abl2rxl] (.clk (\Clks[clk] ), .d (n_200), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[abl2rxl] ));
  CDN_flop \Nanod_reg[rxl2ab] (.clk (\Clks[clk] ), .d (n_201), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[rxl2ab] ));
  CDN_flop \Nanod_reg[rxl2db] (.clk (\Clks[clk] ), .d (n_202), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[rxl2db] ));
  CDN_flop \Nanod_reg[dbh2rxh] (.clk (\Clks[clk] ), .d (n_203), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dbh2rxh] ));
  CDN_flop \Nanod_reg[dbl2rxl] (.clk (\Clks[clk] ), .d (n_204), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[dbl2rxl] ));
  CDN_flop \Nanod_reg[rxh2abh] (.clk (\Clks[clk] ), .d (n_205), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[rxh2abh] ));
  CDN_flop \Nanod_reg[rxh2dbh] (.clk (\Clks[clk] ), .d (n_206), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[rxh2dbh] ));
  CDN_flop \Nanod_reg[isRmc] (.clk (\Clks[clk] ), .d (n_207), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\Nanod[isRmc] ));
  not g170 (n_406, nanoLatch[58]);
  nand g171 (n_407, nanoLatch[57], n_406);
  not g172 (n_116, n_407);
  nand g175 (n_410, nanoLatch[59], n_406);
  not g176 (n_117, n_410);
  nand g179 (n_413, nanoLatch[59], nanoLatch[58]);
  not g180 (n_118, n_413);
  nand g183 (n_416, nanoLatch[58], nanoLatch[57]);
  not g184 (n_119, n_416);
  nand g188 (n_420, nanoLatch[9], n_418, nanoLatch[11]);
  not g5 (n_104, n_420);
  not g191 (n_421, nanoLatch[11]);
  nand g192 (n_424, n_421, nanoLatch[9], nanoLatch[10]);
  not g193 (n_120, n_424);
  nand g197 (n_428, n_425, nanoLatch[10], nanoLatch[11]);
  not g198 (n_121, n_428);
  nand g202 (n_432, n_425, n_418, nanoLatch[11]);
  not g203 (n_122, n_432);
  nor g205 (n_433, nanoLatch[11], nanoLatch[10]);
  nand g206 (n_435, n_433, nanoLatch[9]);
  not g207 (n_103, n_435);
  not g210 (n_436, nanoLatch[31]);
  nand g211 (n_439, n_436, nanoLatch[29], nanoLatch[30]);
  not g212 (n_124, n_439);
  nand g216 (n_443, nanoLatch[29], n_441, nanoLatch[31]);
  not g217 (n_125, n_443);
  nand g221 (n_447, n_444, n_441, nanoLatch[31]);
  not g222 (n_126, n_447);
  nand g226 (n_451, n_436, n_444, nanoLatch[30]);
  not g227 (n_127, n_451);
  nand g230 (n_454, nanoLatch[1], nanoLatch[0]);
  not g231 (n_133, n_454);
  nand g234 (n_457, nanoLatch[1], n_456);
  not g235 (n_160, n_457);
  not g237 (n_459, nanoLatch[1]);
  nand g238 (n_460, nanoLatch[0], n_459);
  not g239 (n_158, n_460);
  nand g242 (n_463, nanoLatch[21], nanoLatch[20]);
  not g243 (\Nanod[au2Pc] , n_463);
  nand g246 (n_466, nanoLatch[21], n_465);
  not g247 (\Nanod[au2Ab] , n_466);
  not g249 (n_468, nanoLatch[21]);
  nand g250 (n_469, nanoLatch[20], n_468);
  not g251 (\Nanod[au2Db] , n_469);
  nand g254 (n_472, nanoLatch[62], n_471);
  not g255 (\Nanod[aluFinish] , n_472);
  not g257 (n_474, nanoLatch[62]);
  nand g258 (n_475, nanoLatch[61], n_474);
  not g259 (\Nanod[aluInit] , n_475);
  nand g262 (n_478, nanoLatch[4], nanoLatch[3]);
  not g263 (\Nanod[au2Aob] , n_478);
  not g265 (n_480, nanoLatch[4]);
  nand g266 (n_481, nanoLatch[3], n_480);
  not g267 (\Nanod[ab2Aob] , n_481);
  nand g270 (n_484, nanoLatch[4], n_483);
  not g271 (\Nanod[db2Aob] , n_484);
  nand g276 (n_489, n_485, n_486, ftuCtrl[1], ftuCtrl[2]);
  not g6 (\Nanod[inl2psw] , n_489);
  nand g281 (n_494, n_486, ftuCtrl[1], ftuCtrl[2], ftuCtrl[3]);
  not g282 (\Nanod[clrTpend] , n_494);
  nand g287 (n_499, ftuCtrl[0], ftuCtrl[1], ftuCtrl[2], ftuCtrl[3]);
  not g288 (n_143, n_499);
  nand g293 (n_504, ftuCtrl[0], ftuCtrl[1], n_502, ftuCtrl[3]);
  not g294 (\Nanod[ssw2Ftu] , n_504);
  nand g299 (n_509, ftuCtrl[0], n_506, n_502, ftuCtrl[3]);
  not g300 (\Nanod[ird2Ftu] , n_509);
  nand g305 (n_514, n_485, ftuCtrl[0], n_506, ftuCtrl[2]);
  not g306 (\Nanod[pswIToFtu] , n_514);
  nand g309 (n_517, nanoLatch[62], nanoLatch[61]);
  not g310 (\Nanod[ftu2Ccr] , n_517);
  nand g315 (n_522, n_485, ftuCtrl[0], ftuCtrl[1], ftuCtrl[2]);
  not g316 (\Nanod[sr2Ftu] , n_522);
  nor g319 (n_525, ftuCtrl[3], ftuCtrl[2]);
  nand g320 (n_526, n_486, ftuCtrl[1], n_525);
  not g321 (\Nanod[ftu2Sr] , n_526);
  nand g326 (n_531, n_486, ftuCtrl[1], n_502, ftuCtrl[3]);
  not g327 (\Nanod[updPren] , n_531);
  nand g332 (n_536, n_486, n_506, ftuCtrl[2], ftuCtrl[3]);
  not g333 (\Nanod[abl2Pren] , n_536);
  nand g338 (n_541, n_486, n_506, n_502, ftuCtrl[3]);
  not g339 (\Nanod[ftu2Abl] , n_541);
  not g343 (n_485, ftuCtrl[3]);
  nand g344 (n_546, n_485, n_486, n_506, ftuCtrl[2]);
  not g345 (n_139, n_546);
  nor g347 (n_547, ftuCtrl[3], ftuCtrl[2], ftuCtrl[1]);
  nand g348 (n_549, n_547, ftuCtrl[0]);
  not g349 (\Nanod[const2Ftu] , n_549);
  nand g354 (n_554, ftuCtrl[0], n_506, ftuCtrl[2], ftuCtrl[3]);
  not g355 (\Nanod[tvn2Ftu] , n_554);
  not g356 (n_418, nanoLatch[10]);
  not g357 (n_486, ftuCtrl[0]);
  not g358 (n_506, ftuCtrl[1]);
  not g359 (n_456, nanoLatch[0]);
  not g360 (n_425, nanoLatch[9]);
  not g361 (n_441, nanoLatch[30]);
  not g362 (n_444, nanoLatch[29]);
  not g363 (n_465, nanoLatch[20]);
  not g364 (n_471, nanoLatch[61]);
  not g365 (n_483, nanoLatch[3]);
  not g366 (n_502, ftuCtrl[2]);
endmodule

module fx68k_and_op_1374(A, Z);
  input [2:0] A;
  output Z;
  wire [2:0] A;
  wire Z;
  wire n_4;
  nand g1 (n_4, A[2], A[1], A[0]);
  not g2 (Z, n_4);
endmodule

module fx68k_or_op_1375(A, Z);
  input [2:0] A;
  output Z;
  wire [2:0] A;
  wire Z;
  wire n_4;
  nor g1 (n_4, A[2], A[1], A[0]);
  not g2 (Z, n_4);
endmodule

module fx68k_and_op_1376(A, Z);
  input [2:0] A;
  output Z;
  wire [2:0] A;
  wire Z;
  wire n_4;
  nand g1 (n_4, A[2], A[1], A[0]);
  not g2 (Z, n_4);
endmodule

module fx68k_equal_unsigned_3572(A, B, Z);
  input [11:0] A, B;
  output Z;
  wire [11:0] A, B;
  wire Z;
  wire n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  xnor g1 (n_26, A[0], B[0]);
  xnor g2 (n_27, A[1], B[1]);
  xnor g3 (n_28, A[2], B[2]);
  xnor g4 (n_29, A[3], B[3]);
  xnor g5 (n_30, A[4], B[4]);
  xnor g6 (n_31, A[5], B[5]);
  xnor g7 (n_32, A[6], B[6]);
  xnor g8 (n_33, A[7], B[7]);
  xnor g9 (n_34, A[8], B[8]);
  xnor g10 (n_35, A[9], B[9]);
  xnor g11 (n_36, A[10], B[10]);
  xnor g12 (n_37, A[11], B[11]);
  nand g13 (n_38, n_26, n_27, n_28, n_29);
  nand g14 (n_39, n_30, n_31, n_32, n_33);
  nand g15 (n_40, n_34, n_35, n_36, n_37);
  nor g16 (Z, n_38, n_39, n_40);
endmodule

module fx68k_bmux_3596(ctl, in_0, in_1, in_2, in_3, z);
  input [1:0] ctl;
  input [3:0] in_0, in_1, in_2, in_3;
  output [3:0] z;
  wire [1:0] ctl;
  wire [3:0] in_0, in_1, in_2, in_3;
  wire [3:0] z;
  CDN_bmux4 g1(.sel0 (ctl[0]), .data0 (in_0[3]), .data1 (in_1[3]),
       .sel1 (ctl[1]), .data2 (in_2[3]), .data3 (in_3[3]), .z (z[3]));
  CDN_bmux4 g2(.sel0 (ctl[0]), .data0 (in_0[2]), .data1 (in_1[2]),
       .sel1 (ctl[1]), .data2 (in_2[2]), .data3 (in_3[2]), .z (z[2]));
  CDN_bmux4 g3(.sel0 (ctl[0]), .data0 (in_0[1]), .data1 (in_1[1]),
       .sel1 (ctl[1]), .data2 (in_2[1]), .data3 (in_3[1]), .z (z[1]));
  CDN_bmux4 g4(.sel0 (ctl[0]), .data0 (in_0[0]), .data1 (in_1[0]),
       .sel1 (ctl[1]), .data2 (in_2[0]), .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_irdDecode(ird, \Irdecod[inhibitCcr] , \Irdecod[macroTvn] ,
     \Irdecod[ftuConst] , \Irdecod[ryIsAreg] , \Irdecod[rxIsAreg] ,
     \Irdecod[ry] , \Irdecod[rx] , \Irdecod[isMovep] , \Irdecod[isByte]
     , \Irdecod[movemPreDecr] , \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp]
     , \Irdecod[ryIsDt] , \Irdecod[rxIsDt] , \Irdecod[toCcr] ,
     \Irdecod[implicitSp] , \Irdecod[isTas] , \Irdecod[isPcRel] );
  input [15:0] ird;
  output \Irdecod[inhibitCcr] , \Irdecod[ryIsAreg] , \Irdecod[rxIsAreg]
       , \Irdecod[isMovep] , \Irdecod[isByte] , \Irdecod[movemPreDecr]
       , \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] ,
       \Irdecod[rxIsDt] , \Irdecod[toCcr] , \Irdecod[implicitSp] ,
       \Irdecod[isTas] , \Irdecod[isPcRel] ;
  output [5:0] \Irdecod[macroTvn] ;
  output [15:0] \Irdecod[ftuConst] ;
  output [2:0] \Irdecod[ry] , \Irdecod[rx] ;
  wire [15:0] ird;
  wire \Irdecod[inhibitCcr] , \Irdecod[ryIsAreg] , \Irdecod[rxIsAreg] ,
       \Irdecod[isMovep] , \Irdecod[isByte] , \Irdecod[movemPreDecr] ,
       \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp] , \Irdecod[ryIsDt] ,
       \Irdecod[rxIsDt] , \Irdecod[toCcr] , \Irdecod[implicitSp] ,
       \Irdecod[isTas] , \Irdecod[isPcRel] ;
  wire [5:0] \Irdecod[macroTvn] ;
  wire [15:0] \Irdecod[ftuConst] ;
  wire [2:0] \Irdecod[ry] , \Irdecod[rx] ;
  wire [15:0] lineOnehot;
  wire [3:0] zero28;
  wire UNCONNECTED483, UNCONNECTED484, eaAreg, eaImmOrAbs, eaIsAreg,
       isDynShift, isRegShift, n_18;
  wire n_26, n_27, n_32, n_33, n_34, n_35, n_36, n_174;
  wire n_175, n_176, n_190, n_191, n_192, n_193, n_194, n_195;
  wire n_198, n_202, n_203, n_204, n_205, n_206, n_208, n_212;
  wire n_214, n_215, n_216, n_217, n_222, n_223, n_225, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_250, n_251, n_256, n_257, n_258, n_259, n_261;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_277, n_278, n_279;
  wire n_281, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_314, n_317, n_319, n_320, n_321, n_322, n_324, n_325;
  wire n_328, n_330, n_334, n_338, n_340, n_345, n_350, n_352;
  wire n_353, n_360, n_363, n_366, n_372, n_404, n_410, n_411;
  wire n_412, n_413, n_414, n_416, n_417, n_418, n_419, n_422;
  wire n_423, n_424, n_425, size11, xIsScc, xStaticMem;
  assign \Irdecod[rx] [0] = ird[9];
  assign \Irdecod[rx] [1] = ird[10];
  assign \Irdecod[rx] [2] = ird[11];
  assign \Irdecod[ry] [0] = ird[0];
  assign \Irdecod[ry] [1] = ird[1];
  assign \Irdecod[ry] [2] = ird[2];
  assign \Irdecod[macroTvn] [4] = 1'b0;
  fx68k_onehotEncoder4 irdLines(ird[15:12], {UNCONNECTED484,
       lineOnehot[14:11], UNCONNECTED483, lineOnehot[9:0]});
  fx68k_and_op_1374 g3(.A (ird[5:3]), .Z (n_243));
  fx68k_or_op_1375 g10(.A (ird[8:6]), .Z (n_204));
  fx68k_and_op_1376 g11(.A (ird[8:6]), .Z (n_205));
  fx68k_equal_unsigned_3572 eq_1059_55(.A (ird[11:0]), .B
       (12'b111001110111), .Z (n_286));
  fx68k_mux_1527 \mux_Irdecod[implicitSp]_1047_10 (.ctl
       ({lineOnehot[6], lineOnehot[4], n_174}), .in_0 (n_175), .in_1
       (n_176), .in_2 (1'b0), .z (\Irdecod[implicitSp] ));
  fx68k_mux_1707 \mux_Irdecod[isByte]_1012_10 (.ctl ({lineOnehot[0],
       lineOnehot[1], lineOnehot[4], lineOnehot[5], n_190, n_191}),
       .in_0 (n_192), .in_1 (1'b1), .in_2 (n_193), .in_3 (n_194), .in_4
       (n_195), .in_5 (1'b0), .z (\Irdecod[isByte] ));
  fx68k_mux_1707 \mux_Irdecod[rxIsAreg]_938_10 (.ctl ({n_198,
       lineOnehot[4], lineOnehot[8], lineOnehot[12], n_202, n_203}),
       .in_0 (n_204), .in_1 (n_205), .in_2 (n_206), .in_3 (n_206),
       .in_4 (n_208), .in_5 (\Irdecod[implicitSp] ), .z
       (\Irdecod[rxIsAreg] ));
  fx68k_mux_1577 \mux_Irdecod[ryIsAreg]_988_10 (.ctl ({lineOnehot[5],
       n_212, lineOnehot[14], n_214}), .in_0 (n_215), .in_1 (1'b0),
       .in_2 (n_216), .in_3 (eaIsAreg), .z (\Irdecod[ryIsAreg] ));
  fx68k_bmux_1504 mux_1066_33(.ctl (n_217), .in_0 ({1'b0, ird[11:9]}),
       .in_1 (4'b1000), .z (zero28));
  fx68k_mux_2286 mux_ftuConst_1069_10(.ctl ({n_212, n_222, n_223,
       lineOnehot[4], n_225}), .in_0 ({ird[7], ird[7], ird[7], ird[7],
       ird[7], ird[7], ird[7], ird[7], ird[7:0]}), .in_1
       ({12'b000000000000, zero28}), .in_2 (16'b0000000000001111),
       .in_3 (16'b0000000010000000), .in_4 (16'b0000000000000000), .z
       (\Irdecod[ftuConst] ));
  fx68k_mux_1527 \mux_Irdecod[macroTvn]_1093_11 (.ctl ({n_234, n_235,
       n_236}), .in_0 (1'b0), .in_1 (1'b0), .in_2 (1'b1), .z (n_241));
  fx68k_bmux_3596 \mux_Irdecod[macroTvn]_1093_65 (.ctl (ird[6:5]),
       .in_0 (4'b0110), .in_1 (4'b0110), .in_2 (ird[3:0]), .in_3
       (4'b0111), .z ({n_240, n_239, n_238, n_237}));
  fx68k_bmux_1854 \mux_Irdecod[macroTvn]_1092_7 (.ctl (lineOnehot[4]),
       .in_0 (5'b00101), .in_1 ({n_241, n_240, n_239, n_238, n_237}),
       .z ({\Irdecod[macroTvn] [5], \Irdecod[macroTvn] [3:0]}));
  and g1 (isRegShift, lineOnehot[14], n_242);
  and g2 (isDynShift, isRegShift, ird[5]);
  and g12 (n_250, eaAreg, ird[8]);
  not g13 (n_251, ird[7]);
  and g14 (n_206, n_250, n_251);
  and g18 (size11, ird[7], ird[6]);
  and g20 (n_256, n_250, n_242);
  or g21 (n_208, size11, n_256);
  not g22 (n_257, ird[8]);
  and g23 (n_258, lineOnehot[4], n_257);
  not g24 (n_259, \Irdecod[implicitSp] );
  and g25 (\Irdecod[rxIsMovem] , n_258, n_259);
  and g27 (n_261, lineOnehot[0], n_257);
  or g28 (\Irdecod[rxIsDt] , lineOnehot[5], n_261);
  not g30 (n_264, ird[1]);
  and g31 (eaImmOrAbs, n_263, n_264);
  not g32 (n_216, isRegShift);
  and g33 (\Irdecod[ryIsDt] , eaImmOrAbs, n_216);
  and g34 (eaIsAreg, n_265, n_266);
  and g35 (n_215, eaIsAreg, n_267);
  and g36 (xIsScc, n_268, n_269);
  and g37 (xStaticMem, n_270, n_271);
  and g38 (n_273, ird[8], n_272);
  and g39 (n_274, n_270, n_272);
  and g41 (n_277, n_275, eaAreg);
  and g44 (n_281, n_278, n_279);
  or g46 (n_193, n_195, \Irdecod[isTas] );
  or g47 (n_194, n_195, xIsScc);
  and g48 (n_283, lineOnehot[0], ird[8]);
  and g49 (\Irdecod[isMovep] , n_283, eaAreg);
  or g50 (n_176, n_284, n_285);
  or g51 (n_288, n_286, n_287);
  and g52 (n_289, lineOnehot[4], n_288);
  and g53 (n_290, lineOnehot[0], n_278);
  or g54 (\Irdecod[toCcr] , n_289, n_290);
  or g56 (n_291, lineOnehot[9], lineOnehot[13]);
  and g57 (n_292, n_291, size11);
  and g58 (n_293, lineOnehot[5], eaAreg);
  or g59 (n_296, n_292, n_293);
  or g60 (n_294, lineOnehot[2], lineOnehot[3]);
  and g61 (n_297, n_294, n_295);
  or g62 (\Irdecod[inhibitCcr] , n_296, n_297);
  not g67 (n_279, xStaticMem);
  nor g69 (n_314, ird[5], ird[4]);
  nand g70 (n_269, n_314, ird[3]);
  not g71 (eaAreg, n_269);
  nand g74 (n_319, n_317, ird[6]);
  not g75 (n_295, n_319);
  nor g77 (n_320, ird[11], ird[10]);
  nand g78 (n_322, n_320, n_321);
  not g79 (n_217, n_322);
  nand g6 (n_328, ird[3], n_324, n_325, ird[6]);
  nor g86 (n_330, n_328, n_251);
  not g87 (n_267, n_330);
  nand g90 (n_242, ird[7], ird[6]);
  nand g93 (n_265, n_314, n_334);
  nor g99 (n_338, ird[11], ird[10], ird[9]);
  nand g100 (n_340, n_338, ird[8]);
  not g101 (n_175, n_340);
  not g107 (n_284, n_345);
  nand g114 (n_353, ird[6], n_251, n_257, n_321);
  nor g116 (n_285, n_352, n_353);
  nand g124 (n_360, n_257, n_321, n_350, ird[11]);
  not g125 (n_270, n_360);
  nand g128 (n_363, ird[8], n_251);
  not g129 (n_275, n_363);
  nor g131 (n_317, ird[8], ird[7]);
  nand g132 (n_366, n_317, n_234);
  not g133 (n_278, n_366);
  not g135 (n_325, ird[5]);
  nand g136 (n_272, n_324, n_325);
  not g137 (n_271, n_272);
  nand g140 (n_372, n_234, n_251);
  not g141 (n_195, n_372);
  nand g149 (n_352, n_350, ird[11]);
  not g154 (n_268, n_242);
  nand g172 (n_345, n_257, ird[9], ird[10], ird[11]);
  nand g177 (n_266, ird[3], ird[4], ird[5]);
  not g178 (n_263, n_266);
  not g184 (n_404, ird[11]);
  nand g185 (n_411, n_404, ird[6], ird[7], n_257);
  nand g186 (n_410, n_321, ird[10]);
  nor g187 (n_287, n_410, n_411);
  not g188 (n_350, ird[10]);
  not g189 (n_334, ird[3]);
  not g190 (n_324, ird[4]);
  not g191 (n_321, ird[9]);
  not g192 (n_234, ird[6]);
  or g193 (n_192, n_273, n_274, n_277, n_281);
  and g194 (n_413, n_412, lineOnehot[4]);
  not g195 (n_412, n_352);
  and g196 (n_414, ird[6], ird[7]);
  and g197 (\Irdecod[isTas] , n_257, ird[9], n_413, n_414);
  and g198 (\Irdecod[movemPreDecr] , \Irdecod[rxIsMovem] , n_334,
       n_324, ird[5]);
  and g199 (n_416, n_284, lineOnehot[4]);
  and g201 (n_417, n_324, ird[5]);
  and g202 (\Irdecod[rxIsUsp] , ird[6], n_251, n_416, n_417);
  and g203 (\Irdecod[isPcRel] , n_418, n_419, n_243, ird[1]);
  not g204 (n_418, isDynShift);
  not g205 (n_419, ird[2]);
  nor g208 (n_174, lineOnehot[4], lineOnehot[6]);
  nor g214 (n_33, lineOnehot[8], lineOnehot[9], lineOnehot[11],
       lineOnehot[12]);
  nor g215 (n_32, lineOnehot[13], lineOnehot[14]);
  nand g216 (n_190, n_32, n_33);
  nor g217 (n_34, lineOnehot[0], lineOnehot[1], lineOnehot[4],
       lineOnehot[5]);
  not g15 (n_35, n_190);
  nand g16 (n_36, n_34, n_35);
  not g17 (n_191, n_36);
  nor g227 (n_422, lineOnehot[1], lineOnehot[2], lineOnehot[3]);
  not g228 (n_198, n_422);
  nor g229 (n_423, lineOnehot[9], lineOnehot[11], lineOnehot[13]);
  not g230 (n_202, n_423);
  nor g231 (n_424, n_198, lineOnehot[4], lineOnehot[8], lineOnehot[12]);
  nand g232 (n_425, n_424, n_423);
  not g233 (n_203, n_425);
  nor g238 (n_18, lineOnehot[7], lineOnehot[6]);
  not g239 (n_212, n_18);
  nor g240 (n_214, lineOnehot[5], n_212, lineOnehot[14]);
  nor g250 (n_26, lineOnehot[14], lineOnehot[5]);
  not g251 (n_222, n_26);
  nor g252 (n_27, lineOnehot[12], lineOnehot[8]);
  not g253 (n_223, n_27);
  nor g254 (n_225, n_212, n_222, n_223, lineOnehot[4]);
  nor g259 (n_235, n_234, n_325);
  nor g261 (n_236, n_234, ird[5]);
endmodule

module fx68k_equal_unsigned_3599(A, B, Z);
  input [31:0] A;
  input [2:0] B;
  output Z;
  wire [31:0] A;
  wire [2:0] B;
  wire Z;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50;
  xnor g1 (n_38, A[0], B[0]);
  xnor g2 (n_39, A[1], B[1]);
  xnor g3 (n_40, A[2], B[2]);
  nor g4 (n_41, A[31], A[30], A[29], A[28]);
  nor g5 (n_42, A[27], A[26], A[25], A[24]);
  nor g6 (n_43, A[23], A[22], A[21], A[20]);
  nor g7 (n_44, A[19], A[18], A[17], A[16]);
  nor g8 (n_45, A[15], A[14], A[13], A[12]);
  nor g9 (n_46, A[11], A[10], A[9], A[8]);
  nor g10 (n_47, A[7], A[6], A[5], A[4]);
  not g11 (n_37, A[3]);
  nand g12 (n_48, n_37, n_38, n_39, n_40);
  nand g13 (n_49, n_41, n_42, n_43, n_44);
  nand g14 (n_50, n_45, n_46, n_47);
  nor g15 (Z, n_48, n_49, n_50);
endmodule

module fx68k_equal_unsigned_3601(A, B, Z);
  input [31:0] A;
  input B;
  output Z;
  wire [31:0] A;
  wire B;
  wire Z;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46;
  xnor g1 (n_35, A[0], B);
  nor g2 (n_36, A[31], A[30], A[29], A[28]);
  nor g3 (n_37, A[27], A[26], A[25], A[24]);
  nor g4 (n_38, A[23], A[22], A[21], A[20]);
  nor g5 (n_39, A[19], A[18], A[17], A[16]);
  nor g6 (n_40, A[15], A[14], A[13], A[12]);
  nor g7 (n_41, A[11], A[10], A[9], A[8]);
  nor g8 (n_42, A[7], A[6], A[5], A[4]);
  nor g9 (n_43, A[3], A[2], A[1]);
  nand g10 (n_45, n_35, n_36, n_37, n_38);
  nand g11 (n_46, n_39, n_40, n_41, n_42);
  not g12 (n_44, n_43);
  nor g13 (Z, n_44, n_45, n_46);
endmodule

module fx68k_equal_unsigned_3603(A, B, Z);
  input [31:0] A;
  input [1:0] B;
  output Z;
  wire [31:0] A;
  wire [1:0] B;
  wire Z;
  wire n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43;
  wire n_44, n_45, n_46, n_47, n_48;
  xnor g1 (n_36, A[0], B[0]);
  xnor g2 (n_37, A[1], B[1]);
  nor g3 (n_38, A[31], A[30], A[29], A[28]);
  nor g4 (n_39, A[27], A[26], A[25], A[24]);
  nor g5 (n_40, A[23], A[22], A[21], A[20]);
  nor g6 (n_41, A[19], A[18], A[17], A[16]);
  nor g7 (n_42, A[15], A[14], A[13], A[12]);
  nor g8 (n_43, A[11], A[10], A[9], A[8]);
  nor g9 (n_44, A[7], A[6], A[5], A[4]);
  nor g10 (n_45, A[3], A[2]);
  nand g11 (n_46, n_36, n_37, n_38, n_39);
  nand g12 (n_47, n_40, n_41, n_42, n_43);
  nand g13 (n_48, n_44, n_45);
  nor g14 (Z, n_46, n_47, n_48);
endmodule

module fx68k_case_box_1412(in_0, out_0);
  input [31:0] in_0;
  output [7:0] out_0;
  wire [31:0] in_0;
  wire [7:0] out_0;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_48, n_63, n_78, n_82, n_83, n_93;
  wire n_108, n_123, n_124, n_125, n_138, n_153, n_166, n_167;
  wire n_168, n_183, n_198, n_208, n_209, n_213, n_228, n_243;
  wire n_250, n_251, n_273, n_274, n_275, n_276, n_288, n_292;
  wire n_293, n_295, n_297, n_299, n_301, n_303, n_305, n_307;
  wire n_309, n_310, n_311, n_318, n_333, n_348, n_363, n_378;
  wire n_393, n_408, n_423, n_489, n_490, n_491, n_492, n_493;
  not g225 (n_273, in_0[31]);
  not g226 (n_274, in_0[30]);
  not g227 (n_33, in_0[29]);
  not g228 (n_48, in_0[28]);
  not g229 (n_63, in_0[27]);
  not g230 (n_78, in_0[26]);
  not g231 (n_93, in_0[25]);
  not g232 (n_108, in_0[24]);
  not g233 (n_123, in_0[23]);
  not g234 (n_138, in_0[22]);
  not g235 (n_153, in_0[21]);
  not g236 (n_168, in_0[20]);
  not g237 (n_183, in_0[19]);
  not g238 (n_198, in_0[18]);
  not g239 (n_213, in_0[17]);
  not g240 (n_228, in_0[16]);
  not g241 (n_243, in_0[15]);
  not g242 (n_275, in_0[14]);
  not g243 (n_276, in_0[13]);
  not g244 (n_288, in_0[12]);
  not g245 (n_303, in_0[11]);
  not g246 (n_318, in_0[10]);
  not g247 (n_333, in_0[9]);
  not g248 (n_348, in_0[8]);
  not g249 (n_363, in_0[7]);
  not g250 (n_378, in_0[6]);
  not g251 (n_393, in_0[5]);
  not g252 (n_408, in_0[4]);
  not g253 (n_423, in_0[3]);
  nand g1 (n_492, n_273, n_274, n_33, n_48);
  nand g2 (n_34, n_63, n_78, n_93, n_108);
  nand g3 (n_35, n_123, n_138, n_153, n_168);
  nand g4 (n_36, n_183, n_198, n_213, n_228);
  nand g5 (n_37, n_243, n_275, n_276, n_288);
  nand g6 (n_38, n_303, n_318, n_333, n_348);
  nand g7 (n_39, n_363, n_378, n_393, n_408);
  nand g8 (n_40, n_423, n_489, n_490, n_491);
  nor g9 (n_42, n_492, n_34, n_35, n_36);
  nor g10 (n_41, n_37, n_38, n_39, n_40);
  nand g11 (n_295, n_41, n_42);
  nand g19 (n_82, n_423, in_0[2], in_0[1], n_491);
  nor g21 (n_83, n_37, n_38, n_39, n_82);
  nand g22 (n_297, n_83, n_42);
  nand g30 (n_124, n_423, n_489, in_0[1], n_491);
  nor g32 (n_125, n_37, n_38, n_39, n_124);
  nand g33 (n_299, n_125, n_42);
  nand g41 (n_166, n_423, n_489, in_0[1], in_0[0]);
  nor g43 (n_167, n_37, n_38, n_39, n_166);
  nand g44 (n_301, n_167, n_42);
  nand g52 (n_208, n_423, in_0[2], n_490, n_491);
  nor g54 (n_209, n_37, n_38, n_39, n_208);
  nand g55 (n_493, n_209, n_42);
  nand g63 (n_250, n_423, in_0[2], n_490, in_0[0]);
  nor g65 (n_251, n_37, n_38, n_39, n_250);
  nand g66 (n_305, n_251, n_42);
  nand g74 (n_292, n_423, n_489, n_490, in_0[0]);
  nor g76 (n_293, n_37, n_38, n_39, n_292);
  nand g77 (n_307, n_293, n_42);
  not g78 (out_0[7], n_295);
  not g79 (out_0[6], n_297);
  not g80 (out_0[5], n_299);
  not g81 (out_0[4], n_301);
  not g82 (out_0[3], n_493);
  not g83 (out_0[2], n_305);
  not g84 (out_0[1], n_307);
  nor g85 (n_310, out_0[7], out_0[6], out_0[5], out_0[4]);
  nor g86 (n_309, out_0[3], out_0[2], out_0[1]);
  nand g87 (n_311, n_309, n_310);
  not g88 (out_0[0], n_311);
  not g89 (n_489, in_0[2]);
  not g90 (n_490, in_0[1]);
  not g91 (n_491, in_0[0]);
endmodule

module fx68k_mux_3623(ctl, in_0, in_1, in_2, in_3, z);
  input [3:0] ctl;
  input [2:0] in_0, in_1, in_2, in_3;
  output [2:0] z;
  wire [3:0] ctl;
  wire [2:0] in_0, in_1, in_2, in_3;
  wire [2:0] z;
  CDN_mux4 g1(.sel0 (ctl[3]), .data0 (in_0[2]), .sel1 (ctl[2]), .data1
       (in_1[2]), .sel2 (ctl[1]), .data2 (in_2[2]), .sel3 (ctl[0]),
       .data3 (in_3[2]), .z (z[2]));
  CDN_mux4 g4(.sel0 (ctl[3]), .data0 (in_0[1]), .sel1 (ctl[2]), .data1
       (in_1[1]), .sel2 (ctl[1]), .data2 (in_2[1]), .sel3 (ctl[0]),
       .data3 (in_3[1]), .z (z[1]));
  CDN_mux4 g5(.sel0 (ctl[3]), .data0 (in_0[0]), .sel1 (ctl[2]), .data1
       (in_1[0]), .sel2 (ctl[1]), .data2 (in_2[0]), .sel3 (ctl[0]),
       .data3 (in_3[0]), .z (z[0]));
endmodule

module fx68k_busControl(\Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] ,
     \Clks[extReset] , \Clks[clk] , enT1, enT4, permStart, permStop,
     iStop, aob0, isWrite, isByte, isRmc, busAvail, bgBlock,
     busAddrErr, waitBusCycle, busStarting, addrOe, bciWrite, rDtack,
     BeDebounced, Vpai, ASn, LDSn, UDSn, eRWn);
  input \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset]
       , \Clks[clk] , enT1, enT4, permStart, permStop, iStop, aob0,
       isWrite, isByte, isRmc, busAvail, rDtack, BeDebounced, Vpai;
  output bgBlock, busAddrErr, waitBusCycle, busStarting, addrOe,
       bciWrite, ASn, LDSn, UDSn, eRWn;
  wire \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset] ,
       \Clks[clk] , enT1, enT4, permStart, permStop, iStop, aob0,
       isWrite, isByte, isRmc, busAvail, rDtack, BeDebounced, Vpai;
  wire bgBlock, busAddrErr, waitBusCycle, busStarting, addrOe,
       bciWrite, ASn, LDSn, UDSn, eRWn;
  wire [31:0] busPhase;
  wire [31:0] next;
  wire UNCONNECTED485, UNCONNECTED486, UNCONNECTED487, UNCONNECTED488,
       UNCONNECTED489, UNCONNECTED490, UNCONNECTED491, UNCONNECTED492;
  wire UNCONNECTED493, UNCONNECTED494, _X_, addrOeDelay, bcComplete,
       bcPend, bcReset, bciByte;
  wire busEnd, busEnding, canStart, isByteT4, isRcmReset, isRmcReg,
       n_5, n_7;
  wire n_8, n_14, n_15, n_16, n_19, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_561, n_562, n_563, n_564;
  wire n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572;
  wire n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580;
  wire n_583, n_586, n_587, n_589, n_590, n_592, n_595, n_596;
  wire n_597, n_598, n_604, n_606, n_607, n_608, n_610, n_613;
  wire n_614, n_615, n_618, n_619, n_620, n_622, n_623, n_624;
  wire n_626, n_629, n_631, n_632, n_634, n_635, n_642, n_643;
  wire n_644, n_645, n_646, n_648, n_649, n_656, n_657, n_658;
  wire n_659, n_660, n_662, n_663, n_664, n_667, n_674, n_675;
  wire n_678, n_680, n_681, n_682, n_683, n_687, n_688, n_884;
  wire n_915, n_923, n_925, n_926, n_927, n_936, rLDS, rUDS;
  wire rmcIdle, wendReg;
  fx68k_equal_unsigned_3599 eq_2314_32(.A (busPhase), .B (3'b101), .Z
       (bcComplete));
  fx68k_equal_unsigned_3601 eq_2302_27(.A (busPhase), .B (1'b1), .Z
       (n_613));
  fx68k_equal_unsigned_3603 eq_2308_33(.A (busPhase), .B (2'b10), .Z
       (busStarting));
  fx68k_equal_unsigned_3599 eq_2328_56(.A (busPhase), .B (3'b110), .Z
       (n_635));
  fx68k_equal_unsigned_3601 eq_2306_25(.A
       ({29'b00000000000000000000000000000, next[2:0]}), .B (1'b1), .Z
       (n_623));
  fx68k_equal_unsigned_3603 eq_2306_43(.A
       ({29'b00000000000000000000000000000, next[2:0]}), .B (2'b10), .Z
       (n_624));
  fx68k_equal_unsigned_3603 eq_2381_50(.A (busPhase), .B (2'b11), .Z
       (n_648));
  fx68k_case_box_1412 ctl_busPhase_2289_9(.in_0 (busPhase), .out_0
       ({n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517}));
  fx68k_mux_1224 mux_next_2289_9(.ctl ({n_510, n_511, n_512, n_513,
       n_514, n_515, n_516, n_517}), .in_0 (5'b00001), .in_1
       (5'b00001), .in_2 (5'b00011), .in_3 (5'b00100), .in_4 ({2'b01,
       _X_, _X_, _X_}), .in_5 ({2'b10, _X_, _X_, _X_}), .in_6 ({2'b11,
       _X_, _X_, _X_}), .in_7 (5'b00001), .z ({n_566, n_565, n_579,
       n_577, n_574}));
  fx68k_bmux_1503 mux_2294_16(.ctl (busEnd), .in_0 (1'b0), .in_1
       (1'b1), .z (n_571));
  fx68k_mux_1577 mux_addrOe_2331_7(.ctl ({\Clks[extReset] , n_523,
       n_524, n_525}), .in_0 (1'b0), .in_1 (1'b1), .in_2 (1'b0), .in_3
       (1'b0), .z (n_656));
  fx68k_bmux_1503 mux_rAS_2367_20(.ctl (n_526), .in_0 (1'b1), .in_1
       (1'b0), .z (n_562));
  fx68k_bmux_1503 mux_rAS_2344_7(.ctl (\Clks[extReset] ), .in_0
       (n_562), .in_1 (1'b1), .z (UNCONNECTED485));
  fx68k_bmux_1520 mux_2295_41(.ctl (canStart), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_564, n_563}));
  fx68k_bmux_1766 mux_2295_16(.ctl (isRcmReset), .in_0 ({1'b0, n_564,
       n_563}), .in_1 (3'b110), .z ({n_578, n_575, n_572}));
  fx68k_bmux_1520 mux_2296_18(.ctl (canStart), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_576, n_573}));
  fx68k_mux_3623 mux_next_2289_87(.ctl ({n_567, n_568, n_569, n_570}),
       .in_0 ({2'b10, n_571}), .in_1 ({n_578, n_575, n_572}), .in_2
       ({1'b0, n_576, n_573}), .in_3 ({n_579, n_577, n_574}), .z
       (next[2:0]));
  fx68k_bmux_1766 mux_busPhase_2282_7(.ctl (\Clks[extReset] ), .in_0
       (next[2:0]), .in_1 (3'b000), .z ({UNCONNECTED488,
       UNCONNECTED487, UNCONNECTED486}));
  fx68k_bmux_1503 mux_wendReg_2419_24(.ctl (n_580), .in_0 (permStop),
       .in_1 (1'b0), .z (n_583));
  fx68k_bmux_1503 mux_wendReg_2411_7(.ctl (\Clks[pwrUp] ), .in_0
       (n_583), .in_1 (1'b0), .z (UNCONNECTED489));
  fx68k_bmux_1503 mux_bciByte_2411_7(.ctl (\Clks[pwrUp] ), .in_0
       (isByteT4), .in_1 (1'b0), .z (UNCONNECTED490));
  fx68k_bmux_1503 mux_isWriteReg_2411_7(.ctl (\Clks[pwrUp] ), .in_0
       (isWrite), .in_1 (1'b0), .z (UNCONNECTED491));
  fx68k_bmux_1503 mux_rRWn_2358_20(.ctl (n_586), .in_0 (1'b0), .in_1
       (1'b1), .z (n_589));
  fx68k_bmux_1503 mux_rRWn_2344_7(.ctl (\Clks[extReset] ), .in_0
       (n_589), .in_1 (1'b1), .z (UNCONNECTED492));
  fx68k_mux_1577 mux_rUDS_2344_7(.ctl ({\Clks[extReset] , n_595, n_596,
       n_597}), .in_0 (1'b1), .in_1 (n_598), .in_2 (n_598), .in_3
       (1'b1), .z (rUDS));
  fx68k_mux_1577 mux_rLDS_2344_7(.ctl ({\Clks[extReset] , n_595, n_596,
       n_597}), .in_0 (1'b1), .in_1 (n_604), .in_2 (n_604), .in_3
       (1'b1), .z (rLDS));
  fx68k_bmux_1503 mux_isRmcReg_2411_7(.ctl (\Clks[pwrUp] ), .in_0
       (n_606), .in_1 (1'b0), .z (UNCONNECTED493));
  fx68k_bmux_1503 mux_bcPend_2419_24(.ctl (n_580), .in_0 (1'b1), .in_1
       (1'b0), .z (n_607));
  fx68k_bmux_1503 mux_bcPend_2411_7(.ctl (\Clks[pwrUp] ), .in_0
       (n_607), .in_1 (1'b0), .z (UNCONNECTED494));
  and g1 (n_608, bcComplete, bcReset);
  and g2 (isRcmReset, n_608, isRmcReg);
  not g3 (n_610, bciByte);
  and g4 (busAddrErr, aob0, n_610);
  not g6 (n_614, ASn);
  and g7 (n_615, n_613, n_614);
  and g8 (rmcIdle, n_615, isRmcReg);
  or g9 (n_618, busAvail, rmcIdle);
  or g10 (n_619, bcPend, permStart);
  and g11 (n_620, n_618, n_619);
  and g14 (canStart, n_620, n_622);
  or g15 (busEnding, n_623, n_624);
  not g16 (n_626, rDtack);
  or g17 (busEnd, n_626, iStop);
  and g19 (n_629, addrOeDelay, BeDebounced);
  and g20 (n_631, n_629, Vpai);
  or g21 (bcReset, \Clks[extReset] , n_631);
  and g23 (waitBusCycle, wendReg, n_632);
  and g24 (n_634, busStarting, ASn);
  or g25 (bgBlock, n_634, n_635);
  and g26 (n_7, \Clks[enPhi2] , busStarting);
  and g27 (n_8, \Clks[enPhi1] , n_635);
  not g28 (n_561, isRmcReg);
  and g31 (n_586, \Clks[enPhi1] , busEnding);
  and g32 (n_587, \Clks[enPhi1] , bciWrite);
  and g34 (n_526, \Clks[enPhi1] , busStarting);
  and g35 (n_527, \Clks[enPhi2] , n_635);
  and g36 (n_528, \Clks[enPhi2] , bcComplete);
  not g40 (n_642, bciWrite);
  and g42 (n_590, n_642, n_643);
  not g43 (n_644, aob0);
  or g44 (n_645, n_610, n_644);
  not g45 (n_598, n_645);
  or g46 (n_646, n_610, aob0);
  not g47 (n_604, n_646);
  and g49 (n_649, n_587, n_648);
  and g51 (n_592, n_649, n_643);
  or g65 (n_678, bcComplete, bcReset);
  and g66 (n_580, \Clks[enPhi2] , n_678);
  and g67 (n_518, enT1, permStart);
  not g68 (n_680, isWrite);
  and g69 (n_606, isRmc, n_680);
  CDN_dc logicX_inst(.cf (1'b0), .dcf (1'b1), .z (_X_));
  not g76 (n_15, \Clks[extReset] );
  not g82 (n_659, n_527);
  not g88 (n_681, n_580);
  and g99 (n_658, n_561, n_528);
  and g100 (n_660, n_658, n_659);
  or g101 (n_662, n_660, n_527);
  and g102 (n_663, n_526, n_15);
  and g103 (n_664, n_590, n_595);
  or g113 (n_675, n_674, n_586);
  and g114 (n_682, n_518, n_681);
  or g115 (n_683, n_682, n_580);
  and g119 (n_687, enT1, n_681);
  or g120 (n_688, n_687, n_580);
  CDN_flop \busPhase_reg[0] (.clk (\Clks[clk] ), .d (next[0]), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[0]));
  CDN_flop \busPhase_reg[1] (.clk (\Clks[clk] ), .d (next[1]), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[1]));
  CDN_flop \busPhase_reg[2] (.clk (\Clks[clk] ), .d (next[2]), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[2]));
  CDN_flop \busPhase_reg[3] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[3]));
  CDN_flop \busPhase_reg[4] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[4]));
  CDN_flop \busPhase_reg[5] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[5]));
  CDN_flop \busPhase_reg[6] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[6]));
  CDN_flop \busPhase_reg[7] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[7]));
  CDN_flop \busPhase_reg[8] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[8]));
  CDN_flop \busPhase_reg[9] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[9]));
  CDN_flop \busPhase_reg[10] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[10]));
  CDN_flop \busPhase_reg[11] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[11]));
  CDN_flop \busPhase_reg[12] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[12]));
  CDN_flop \busPhase_reg[13] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[13]));
  CDN_flop \busPhase_reg[14] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[14]));
  CDN_flop \busPhase_reg[15] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[15]));
  CDN_flop \busPhase_reg[16] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[16]));
  CDN_flop \busPhase_reg[17] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[17]));
  CDN_flop \busPhase_reg[18] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[18]));
  CDN_flop \busPhase_reg[19] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[19]));
  CDN_flop \busPhase_reg[20] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[20]));
  CDN_flop \busPhase_reg[21] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[21]));
  CDN_flop \busPhase_reg[22] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[22]));
  CDN_flop \busPhase_reg[23] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[23]));
  CDN_flop \busPhase_reg[24] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[24]));
  CDN_flop \busPhase_reg[25] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[25]));
  CDN_flop \busPhase_reg[26] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[26]));
  CDN_flop \busPhase_reg[27] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[27]));
  CDN_flop \busPhase_reg[28] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[28]));
  CDN_flop \busPhase_reg[29] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[29]));
  CDN_flop \busPhase_reg[30] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[30]));
  CDN_flop \busPhase_reg[31] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (busPhase[31]));
  not g184 (n_622, bcReset);
  not g185 (n_632, bcComplete);
  not g216 (n_643, busAddrErr);
  CDN_flop addrOe_reg(.clk (\Clks[clk] ), .d (n_656), .sena (n_657),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (addrOe));
  CDN_flop rAS_reg(.clk (\Clks[clk] ), .d (1'b1), .sena (n_662), .aclr
       (1'b0), .apre (1'b0), .srl (n_884), .srd (\Clks[extReset] ), .q
       (ASn));
  or g219 (n_884, n_663, \Clks[extReset] );
  CDN_flop rLDS_reg(.clk (\Clks[clk] ), .d (rLDS), .sena (n_667), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (LDSn));
  CDN_flop rUDS_reg(.clk (\Clks[clk] ), .d (rUDS), .sena (n_667), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (UDSn));
  CDN_flop rRWn_reg(.clk (\Clks[clk] ), .d (n_589), .sena (n_675),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b1), .q (eRWn));
  CDN_flop addrOeDelay_reg(.clk (\Clks[clk] ), .d (addrOe), .sena
       (\Clks[enPhi1] ), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (addrOeDelay));
  CDN_flop isByteT4_reg(.clk (\Clks[clk] ), .d (isByte), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (isByteT4));
  CDN_flop bcPend_reg(.clk (\Clks[clk] ), .d (n_607), .sena (n_683),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd (1'b0),
       .q (bcPend));
  CDN_flop isWriteReg_reg(.clk (\Clks[clk] ), .d (isWrite), .sena
       (n_682), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (bciWrite));
  CDN_flop bciByte_reg(.clk (\Clks[clk] ), .d (isByteT4), .sena
       (n_682), .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd
       (1'b0), .q (bciByte));
  CDN_flop isRmcReg_reg(.clk (\Clks[clk] ), .d (n_606), .sena (n_682),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd (1'b0),
       .q (isRmcReg));
  CDN_flop wendReg_reg(.clk (\Clks[clk] ), .d (n_583), .sena (n_688),
       .aclr (1'b0), .apre (1'b0), .srl (\Clks[pwrUp] ), .srd (1'b0),
       .q (wendReg));
  or g238 (n_657, n_525, n_524, n_523, \Clks[extReset] );
  or g239 (n_667, n_597, n_596, n_664, \Clks[extReset] );
  and g241 (n_674, n_915, busStarting, bciWrite, n_587);
  not g242 (n_915, n_586);
  or g243 (n_14, n_7, \Clks[extReset] );
  and g246 (n_523, n_15, n_7);
  not g5 (n_16, n_14);
  and g247 (n_524, n_16, n_8);
  nor g255 (n_567, n_19, n_566);
  not g256 (n_19, n_565);
  nor g257 (n_568, n_565, n_5);
  not g258 (n_5, n_566);
  nor g259 (n_569, n_19, n_5);
  nor g260 (n_570, n_565, n_566);
  or g273 (n_923, n_526, \Clks[extReset] );
  or g274 (n_926, n_592, n_923);
  and g276 (n_595, n_15, n_526);
  not g277 (n_925, n_923);
  and g278 (n_596, n_925, n_592);
  not g279 (n_927, n_926);
  and g280 (n_597, n_927, n_528);
  nor g285 (n_936, n_8, n_14);
  and g286 (n_525, \Clks[enPhi1] , n_561, busEnding, n_936);
endmodule

module fx68k_case_box_1428(in_0, out_0);
  input [31:0] in_0;
  output [8:0] out_0;
  wire [31:0] in_0;
  wire [8:0] out_0;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_54, n_71, n_82, n_83, n_88, n_105;
  wire n_122, n_124, n_125, n_139, n_156, n_166, n_167, n_173;
  wire n_190, n_207, n_208, n_209, n_224, n_241, n_250, n_251;
  wire n_258, n_275, n_307, n_308, n_309, n_310, n_326, n_334;
  wire n_335, n_337, n_339, n_341, n_343, n_345, n_347, n_349;
  wire n_351, n_353, n_354, n_355, n_360, n_377, n_394, n_411;
  wire n_428, n_445, n_462, n_479, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560;
  not g257 (n_307, in_0[31]);
  not g258 (n_308, in_0[30]);
  not g259 (n_37, in_0[29]);
  not g260 (n_54, in_0[28]);
  not g261 (n_71, in_0[27]);
  not g262 (n_88, in_0[26]);
  not g263 (n_105, in_0[25]);
  not g264 (n_122, in_0[24]);
  not g265 (n_139, in_0[23]);
  not g266 (n_156, in_0[22]);
  not g267 (n_173, in_0[21]);
  not g268 (n_190, in_0[20]);
  not g269 (n_207, in_0[19]);
  not g270 (n_224, in_0[18]);
  not g271 (n_241, in_0[17]);
  not g272 (n_258, in_0[16]);
  not g273 (n_275, in_0[15]);
  not g274 (n_309, in_0[14]);
  not g275 (n_310, in_0[13]);
  not g276 (n_326, in_0[12]);
  not g277 (n_343, in_0[11]);
  not g278 (n_360, in_0[10]);
  not g279 (n_377, in_0[9]);
  not g280 (n_394, in_0[8]);
  not g281 (n_411, in_0[7]);
  not g282 (n_428, in_0[6]);
  not g283 (n_445, in_0[5]);
  not g284 (n_462, in_0[4]);
  not g285 (n_479, in_0[3]);
  nand g1 (n_33, n_307, n_308, n_37, n_54);
  nand g2 (n_34, n_71, n_88, n_105, n_122);
  nand g3 (n_35, n_139, n_156, n_173, n_190);
  nand g4 (n_36, n_207, n_224, n_241, n_258);
  nand g5 (n_557, n_275, n_309, n_310, n_326);
  nand g6 (n_38, n_343, n_360, n_377, n_394);
  nand g7 (n_39, n_411, n_428, n_445, n_462);
  nand g8 (n_40, n_479, n_554, n_555, n_556);
  nor g9 (n_42, n_33, n_34, n_35, n_36);
  nor g10 (n_41, n_557, n_38, n_39, n_40);
  nand g11 (n_337, n_41, n_42);
  nand g19 (n_82, n_479, n_554, n_555, in_0[0]);
  nor g21 (n_83, n_557, n_38, n_39, n_82);
  nand g22 (n_339, n_83, n_42);
  nand g30 (n_124, n_479, in_0[2], n_555, n_556);
  nor g32 (n_125, n_557, n_38, n_39, n_124);
  nand g33 (n_341, n_125, n_42);
  nand g41 (n_166, n_479, n_554, in_0[1], n_556);
  nor g43 (n_167, n_557, n_38, n_39, n_166);
  nand g44 (n_560, n_167, n_42);
  nand g52 (n_208, n_479, n_554, in_0[1], in_0[0]);
  nor g54 (n_209, n_557, n_38, n_39, n_208);
  nand g55 (n_345, n_209, n_42);
  nand g63 (n_250, n_479, in_0[2], in_0[1], n_556);
  nor g65 (n_251, n_557, n_38, n_39, n_250);
  nand g66 (n_347, n_251, n_42);
  nand g74 (n_558, n_479, in_0[2], n_555, in_0[0]);
  nor g76 (n_559, n_557, n_38, n_39, n_558);
  nand g77 (n_349, n_559, n_42);
  nand g85 (n_334, n_479, in_0[2], in_0[1], in_0[0]);
  nor g87 (n_335, n_557, n_38, n_39, n_334);
  nand g88 (n_351, n_335, n_42);
  not g89 (out_0[8], n_337);
  not g90 (out_0[7], n_339);
  not g91 (out_0[6], n_341);
  not g92 (out_0[5], n_560);
  not g93 (out_0[4], n_345);
  not g94 (out_0[3], n_347);
  not g95 (out_0[2], n_349);
  not g96 (out_0[1], n_351);
  nor g97 (n_354, out_0[8], out_0[7], out_0[6], out_0[5]);
  nor g98 (n_353, out_0[4], out_0[3], out_0[2], out_0[1]);
  nand g99 (n_355, n_353, n_354);
  not g100 (out_0[0], n_355);
  not g101 (n_554, in_0[2]);
  not g102 (n_555, in_0[1]);
  not g103 (n_556, in_0[0]);
endmodule

module fx68k_mux_3637(ctl, in_0, in_1, in_2, in_3, in_4, in_5, in_6,
     in_7, in_8, z);
  input [8:0] ctl;
  input [5:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  output [5:0] z;
  wire [8:0] ctl;
  wire [5:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8;
  wire [5:0] z;
  CDN_mux9 g1(.sel0 (ctl[8]), .data0 (in_0[5]), .sel1 (ctl[7]), .data1
       (in_1[5]), .sel2 (ctl[6]), .data2 (in_2[5]), .sel3 (ctl[5]),
       .data3 (in_3[5]), .sel4 (ctl[4]), .data4 (in_4[5]), .sel5
       (ctl[3]), .data5 (in_5[5]), .sel6 (ctl[2]), .data6 (in_6[5]),
       .sel7 (ctl[1]), .data7 (in_7[5]), .sel8 (ctl[0]), .data8
       (in_8[5]), .z (z[5]));
  CDN_mux9 g7(.sel0 (ctl[8]), .data0 (in_0[4]), .sel1 (ctl[7]), .data1
       (in_1[4]), .sel2 (ctl[6]), .data2 (in_2[4]), .sel3 (ctl[5]),
       .data3 (in_3[4]), .sel4 (ctl[4]), .data4 (in_4[4]), .sel5
       (ctl[3]), .data5 (in_5[4]), .sel6 (ctl[2]), .data6 (in_6[4]),
       .sel7 (ctl[1]), .data7 (in_7[4]), .sel8 (ctl[0]), .data8
       (in_8[4]), .z (z[4]));
  CDN_mux9 g8(.sel0 (ctl[8]), .data0 (in_0[3]), .sel1 (ctl[7]), .data1
       (in_1[3]), .sel2 (ctl[6]), .data2 (in_2[3]), .sel3 (ctl[5]),
       .data3 (in_3[3]), .sel4 (ctl[4]), .data4 (in_4[3]), .sel5
       (ctl[3]), .data5 (in_5[3]), .sel6 (ctl[2]), .data6 (in_6[3]),
       .sel7 (ctl[1]), .data7 (in_7[3]), .sel8 (ctl[0]), .data8
       (in_8[3]), .z (z[3]));
  CDN_mux9 g9(.sel0 (ctl[8]), .data0 (in_0[2]), .sel1 (ctl[7]), .data1
       (in_1[2]), .sel2 (ctl[6]), .data2 (in_2[2]), .sel3 (ctl[5]),
       .data3 (in_3[2]), .sel4 (ctl[4]), .data4 (in_4[2]), .sel5
       (ctl[3]), .data5 (in_5[2]), .sel6 (ctl[2]), .data6 (in_6[2]),
       .sel7 (ctl[1]), .data7 (in_7[2]), .sel8 (ctl[0]), .data8
       (in_8[2]), .z (z[2]));
  CDN_mux9 g10(.sel0 (ctl[8]), .data0 (in_0[1]), .sel1 (ctl[7]), .data1
       (in_1[1]), .sel2 (ctl[6]), .data2 (in_2[1]), .sel3 (ctl[5]),
       .data3 (in_3[1]), .sel4 (ctl[4]), .data4 (in_4[1]), .sel5
       (ctl[3]), .data5 (in_5[1]), .sel6 (ctl[2]), .data6 (in_6[1]),
       .sel7 (ctl[1]), .data7 (in_7[1]), .sel8 (ctl[0]), .data8
       (in_8[1]), .z (z[1]));
  CDN_mux9 g11(.sel0 (ctl[8]), .data0 (in_0[0]), .sel1 (ctl[7]), .data1
       (in_1[0]), .sel2 (ctl[6]), .data2 (in_2[0]), .sel3 (ctl[5]),
       .data3 (in_3[0]), .sel4 (ctl[4]), .data4 (in_4[0]), .sel5
       (ctl[3]), .data5 (in_5[0]), .sel6 (ctl[2]), .data6 (in_6[0]),
       .sel7 (ctl[1]), .data7 (in_7[0]), .sel8 (ctl[0]), .data8
       (in_8[0]), .z (z[0]));
endmodule

module fx68k_case_box_1429(in_0, out_0);
  input [1:0] in_0;
  output [3:0] out_0;
  wire [1:0] in_0;
  wire [3:0] out_0;
  wire n_3, n_6, n_9, n_15, n_23, n_24;
  nand g1 (n_9, in_0[0], in_0[1]);
  nand g2 (n_23, n_3, in_0[1]);
  nand g3 (n_24, in_0[0], n_6);
  nand g4 (n_15, n_3, n_6);
  not g5 (out_0[3], n_9);
  not g6 (out_0[2], n_23);
  not g7 (out_0[1], n_24);
  not g8 (out_0[0], n_15);
  not g11 (n_3, in_0[0]);
  not g12 (n_6, in_0[1]);
endmodule

module fx68k_mux_3649(ctl, in_0, in_1, in_2, in_3, in_4, z);
  input [4:0] ctl;
  input [2:0] in_0, in_1, in_2, in_3, in_4;
  output [2:0] z;
  wire [4:0] ctl;
  wire [2:0] in_0, in_1, in_2, in_3, in_4;
  wire [2:0] z;
  CDN_mux5 g1(.sel0 (ctl[4]), .data0 (in_0[2]), .sel1 (ctl[3]), .data1
       (in_1[2]), .sel2 (ctl[2]), .data2 (in_2[2]), .sel3 (ctl[1]),
       .data3 (in_3[2]), .sel4 (ctl[0]), .data4 (in_4[2]), .z (z[2]));
  CDN_mux5 g4(.sel0 (ctl[4]), .data0 (in_0[1]), .sel1 (ctl[3]), .data1
       (in_1[1]), .sel2 (ctl[2]), .data2 (in_2[1]), .sel3 (ctl[1]),
       .data3 (in_3[1]), .sel4 (ctl[0]), .data4 (in_4[1]), .z (z[1]));
  CDN_mux5 g5(.sel0 (ctl[4]), .data0 (in_0[0]), .sel1 (ctl[3]), .data1
       (in_1[0]), .sel2 (ctl[2]), .data2 (in_2[0]), .sel3 (ctl[1]),
       .data3 (in_3[0]), .sel4 (ctl[0]), .data4 (in_4[0]), .z (z[0]));
endmodule

module fx68k_case_box_1435(in_0, out_0);
  input [31:0] in_0;
  output [1:0] out_0;
  wire [31:0] in_0;
  wire [1:0] out_0;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_48, n_57, n_66, n_75, n_82, n_83;
  wire n_84, n_93, n_102, n_111, n_120, n_124, n_125, n_129;
  wire n_138, n_147, n_156, n_157, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_174, n_183, n_192, n_201;
  wire n_210, n_219, n_228, n_237, n_246, n_255, n_291, n_292;
  wire n_293, n_294, n_295, n_296;
  not g1 (out_0[0], out_0[1]);
  not g129 (n_165, in_0[31]);
  not g130 (n_166, in_0[30]);
  not g131 (n_167, in_0[29]);
  not g132 (n_168, in_0[28]);
  not g133 (n_39, in_0[27]);
  not g134 (n_48, in_0[26]);
  not g135 (n_57, in_0[25]);
  not g136 (n_66, in_0[24]);
  not g137 (n_75, in_0[23]);
  not g138 (n_84, in_0[22]);
  not g139 (n_93, in_0[21]);
  not g140 (n_102, in_0[20]);
  not g141 (n_111, in_0[19]);
  not g142 (n_120, in_0[18]);
  not g143 (n_129, in_0[17]);
  not g144 (n_138, in_0[16]);
  not g145 (n_147, in_0[15]);
  not g146 (n_156, in_0[14]);
  not g147 (n_169, in_0[13]);
  not g148 (n_174, in_0[12]);
  not g149 (n_183, in_0[11]);
  not g150 (n_192, in_0[10]);
  not g151 (n_201, in_0[9]);
  not g152 (n_210, in_0[8]);
  not g153 (n_219, in_0[7]);
  not g154 (n_228, in_0[6]);
  not g155 (n_237, in_0[5]);
  not g156 (n_246, in_0[4]);
  not g157 (n_255, in_0[3]);
  nand g162 (n_33, n_165, n_166, n_167, n_168);
  nand g2 (n_34, n_39, n_48, n_57, n_66);
  nand g3 (n_35, n_75, n_84, n_93, n_102);
  nand g4 (n_36, n_111, n_120, n_129, n_138);
  nand g5 (n_37, n_147, n_156, n_169, n_174);
  nand g6 (n_38, n_183, n_192, n_201, n_210);
  nand g7 (n_293, n_219, n_228, n_237, n_246);
  nand g8 (n_40, n_255, n_291, in_0[1], n_292);
  nor g9 (n_42, n_33, n_34, n_35, n_36);
  nor g10 (n_41, n_37, n_38, n_293, n_40);
  nand g11 (n_296, n_41, n_42);
  nand g19 (n_82, n_255, in_0[2], in_0[1], n_292);
  nor g21 (n_83, n_37, n_38, n_293, n_82);
  nand g22 (n_170, n_83, n_42);
  nand g30 (n_124, n_255, n_291, in_0[1], in_0[0]);
  nor g32 (n_125, n_37, n_38, n_293, n_124);
  nand g33 (n_171, n_125, n_42);
  nand g41 (n_294, n_255, in_0[2], n_157, in_0[0]);
  nor g43 (n_295, n_37, n_38, n_293, n_294);
  nand g44 (n_172, n_295, n_42);
  nand g45 (out_0[1], n_296, n_170, n_171, n_172);
  not g47 (n_291, in_0[2]);
  not g48 (n_292, in_0[0]);
  not g49 (n_157, in_0[1]);
endmodule

module fx68k_busArbiter(\Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] ,
     \Clks[extReset] , \Clks[clk] , BRi, BgackI, Halti, bgBlock,
     busAvail, BGn);
  input \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset]
       , \Clks[clk] , BRi, BgackI, Halti, bgBlock;
  output busAvail, BGn;
  wire \Clks[enPhi2] , \Clks[enPhi1] , \Clks[pwrUp] , \Clks[extReset] ,
       \Clks[clk] , BRi, BgackI, Halti, bgBlock;
  wire busAvail, BGn;
  wire [31:0] dmaPhase;
  wire [31:0] next;
  wire UNCONNECTED495, UNCONNECTED496, UNCONNECTED497, UNCONNECTED498,
       UNCONNECTED499, _X_, granting, n_6;
  wire n_13, n_15, n_33, n_34, n_35, n_36, n_642, n_643;
  wire n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_652;
  wire n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660;
  wire n_661, n_662, n_663, n_666, n_667, n_668, n_669, n_670;
  wire n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678;
  wire n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686;
  wire n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_695;
  wire n_697, rGranted;
  fx68k_case_box_1428 ctl_dmaPhase_2163_8(.in_0 (dmaPhase), .out_0
       ({n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649,
       n_650}));
  fx68k_mux_3637 mux_next_2163_8(.ctl ({n_642, n_643, n_644, n_645,
       n_646, n_647, n_648, n_649, n_650}), .in_0 (6'b000001), .in_1
       ({3'b001, _X_, _X_, _X_}), .in_2 ({3'b010, _X_, _X_, _X_}),
       .in_3 (6'b000011), .in_4 ({3'b011, _X_, _X_, _X_}), .in_5
       (6'b000101), .in_6 ({3'b100, _X_, _X_, _X_}), .in_7 (6'b000100),
       .in_8 (6'b000001), .z ({n_672, n_671, n_670, n_691, n_686,
       n_681}));
  fx68k_bmux_1520 mux_next_2170_14(.ctl (n_653), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_655, n_654}));
  fx68k_bmux_1766 mux_next_2168_14(.ctl (n_652), .in_0 ({1'b0, n_655,
       n_654}), .in_1 (3'b100), .z ({n_658, n_657, n_656}));
  fx68k_bmux_1766 mux_next_2166_9(.ctl (bgBlock), .in_0 ({n_658, n_657,
       n_656}), .in_1 (3'b001), .z ({n_687, n_682, n_678}));
  fx68k_bmux_1520 mux_next_2179_22(.ctl (n_660), .in_0 (2'b01), .in_1
       (2'b10), .z ({n_662, n_661}));
  fx68k_bmux_1766 mux_next_2177_14(.ctl (n_659), .in_0 ({n_662, 1'b0,
       n_661}), .in_1 (3'b110), .z ({n_688, n_683, n_679}));
  fx68k_bmux_1766 mux_2186_21(.ctl (n_663), .in_0 (3'b100), .in_1
       (3'b011), .z ({n_689, n_684, n_680}));
  fx68k_case_box_1429 ctl_2190_5(.in_0 ({BgackI, BRi}), .out_0 ({n_666,
       n_667, n_668, n_669}));
  fx68k_mux_1696 mux_next_2190_5(.ctl ({n_666, n_667, n_668, n_669}),
       .in_0 (2'b00), .in_1 (2'b01), .in_2 (2'b11), .in_3 (2'b10), .z
       ({n_690, n_685}));
  fx68k_mux_3649 mux_next_2163_25(.ctl ({n_673, n_674, n_675, n_676,
       n_677}), .in_0 ({n_687, n_682, n_678}), .in_1 ({n_688, n_683,
       n_679}), .in_2 ({n_689, n_684, n_680}), .in_3 ({n_690, n_685,
       1'b1}), .in_4 ({n_691, n_686, n_681}), .z (next[2:0]));
  fx68k_case_box_1435 ctl_next_2209_16(.in_0
       ({29'b00000000000000000000000000000, next[2:0]}), .out_0
       ({n_692, n_693}));
  fx68k_mux_1783 mux_granting_2209_16(.ctl ({n_692, n_693}), .in_0
       (1'b1), .in_1 (1'b0), .z (granting));
  fx68k_bmux_1503 mux_rGranted_2219_7(.ctl (\Clks[extReset] ), .in_0
       (granting), .in_1 (1'b0), .z (UNCONNECTED495));
  fx68k_bmux_1503 mux_BGn_2230_7(.ctl (\Clks[extReset] ), .in_0
       (n_695), .in_1 (1'b1), .z (UNCONNECTED496));
  fx68k_bmux_1766 mux_dmaPhase_2219_7(.ctl (\Clks[extReset] ), .in_0
       (next[2:0]), .in_1 (3'b000), .z ({UNCONNECTED499,
       UNCONNECTED498, UNCONNECTED497}));
  not g1 (n_652, BgackI);
  not g2 (n_653, BRi);
  and g5 (n_659, n_653, n_697);
  and g7 (n_660, n_652, n_697);
  and g9 (n_663, n_653, BgackI);
  not g12 (n_695, rGranted);
  CDN_dc logicX_inst(.cf (1'b0), .dcf (1'b1), .z (_X_));
  not g27 (n_697, bgBlock);
  CDN_flop BGn_reg(.clk (\Clks[clk] ), .d (n_695), .sena (\Clks[enPhi1]
       ), .aclr (1'b0), .apre (1'b0), .srl (\Clks[extReset] ), .srd
       (1'b1), .q (BGn));
  CDN_flop \dmaPhase_reg[0] (.clk (\Clks[clk] ), .d (next[0]), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[0]));
  CDN_flop \dmaPhase_reg[1] (.clk (\Clks[clk] ), .d (next[1]), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[1]));
  CDN_flop \dmaPhase_reg[2] (.clk (\Clks[clk] ), .d (next[2]), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[2]));
  CDN_flop \dmaPhase_reg[3] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[3]));
  CDN_flop \dmaPhase_reg[4] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[4]));
  CDN_flop \dmaPhase_reg[5] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[5]));
  CDN_flop \dmaPhase_reg[6] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[6]));
  CDN_flop \dmaPhase_reg[7] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[7]));
  CDN_flop \dmaPhase_reg[8] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[8]));
  CDN_flop \dmaPhase_reg[9] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[9]));
  CDN_flop \dmaPhase_reg[10] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[10]));
  CDN_flop \dmaPhase_reg[11] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[11]));
  CDN_flop \dmaPhase_reg[12] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[12]));
  CDN_flop \dmaPhase_reg[13] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[13]));
  CDN_flop \dmaPhase_reg[14] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[14]));
  CDN_flop \dmaPhase_reg[15] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[15]));
  CDN_flop \dmaPhase_reg[16] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[16]));
  CDN_flop \dmaPhase_reg[17] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[17]));
  CDN_flop \dmaPhase_reg[18] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[18]));
  CDN_flop \dmaPhase_reg[19] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[19]));
  CDN_flop \dmaPhase_reg[20] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[20]));
  CDN_flop \dmaPhase_reg[21] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[21]));
  CDN_flop \dmaPhase_reg[22] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[22]));
  CDN_flop \dmaPhase_reg[23] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[23]));
  CDN_flop \dmaPhase_reg[24] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[24]));
  CDN_flop \dmaPhase_reg[25] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[25]));
  CDN_flop \dmaPhase_reg[26] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[26]));
  CDN_flop \dmaPhase_reg[27] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[27]));
  CDN_flop \dmaPhase_reg[28] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[28]));
  CDN_flop \dmaPhase_reg[29] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[29]));
  CDN_flop \dmaPhase_reg[30] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[30]));
  CDN_flop \dmaPhase_reg[31] (.clk (\Clks[clk] ), .d (1'b0), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (dmaPhase[31]));
  CDN_flop rGranted_reg(.clk (\Clks[clk] ), .d (granting), .sena
       (\Clks[enPhi2] ), .aclr (1'b0), .apre (1'b0), .srl
       (\Clks[extReset] ), .srd (1'b0), .q (rGranted));
  and g92 (busAvail, Halti, BRi, BgackI, n_695);
  nand g93 (n_13, n_33, n_34, n_670);
  nand g94 (n_15, n_33, n_671, n_6);
  nand g3 (n_35, n_33, n_671, n_670);
  nand g4 (n_36, n_672, n_34, n_6);
  not g95 (n_673, n_13);
  not g6 (n_674, n_15);
  not g96 (n_675, n_35);
  not g8 (n_676, n_36);
  nor g97 (n_677, n_673, n_674, n_675, n_676);
  not g10 (n_33, n_672);
  not g11 (n_34, n_671);
  not g98 (n_6, n_670);
endmodule

module fx68k_not_op_1441(A, Z);
  input [2:0] A;
  output [2:0] Z;
  wire [2:0] A;
  wire [2:0] Z;
  not g1 (Z[2], A[2]);
  not g2 (Z[1], A[1]);
  not g3 (Z[0], A[0]);
endmodule

module fx68k_gt_unsigned(A, B, Z);
  input [2:0] A, B;
  output Z;
  wire [2:0] A, B;
  wire Z;
  wire n_13, n_14, n_16, n_17, n_19, n_20, n_21, n_22;
  wire n_23, n_24, n_25, n_26, n_27, n_28;
  not g2 (n_13, A[2]);
  not g3 (n_14, A[1]);
  not g5 (Z, n_16);
  nand g9 (n_20, n_17, A[0]);
  nor g10 (n_19, B[1], n_14);
  nand g11 (n_22, B[1], n_14);
  nor g12 (n_24, B[2], n_13);
  nand g13 (n_27, B[2], n_13);
  not g14 (n_21, n_19);
  nand g15 (n_23, n_20, n_21);
  nand g16 (n_25, n_22, n_23);
  not g17 (n_26, n_24);
  nand g18 (n_28, n_25, n_26);
  nand g19 (n_16, n_27, n_28);
  not g25 (n_17, B[0]);
endmodule

module fx68k_add_unsigned_3681(A, B, Z);
  input [3:0] A;
  input B;
  output [3:0] Z;
  wire [3:0] A;
  wire B;
  wire [3:0] Z;
  wire n_11, n_18, n_21, n_28, n_30, n_34, n_35, n_37;
  wire n_38;
  xor g1 (Z[0], A[0], B);
  nand g2 (n_11, A[0], B);
  nand g13 (n_21, n_18, A[1]);
  nand g20 (n_30, n_28, A[2]);
  xnor g25 (Z[1], n_18, n_34);
  xnor g27 (Z[2], n_28, n_35);
  xnor g30 (Z[3], n_37, n_38);
  not g35 (n_18, n_11);
  not g36 (n_34, A[1]);
  not g37 (n_35, A[2]);
  not g38 (n_38, A[3]);
  not g39 (n_28, n_21);
  not g40 (n_37, n_30);
endmodule

module fx68k_bmux_3758(ctl, in_0, in_1, z);
  input ctl;
  input [67:0] in_0, in_1;
  output [67:0] z;
  wire ctl;
  wire [67:0] in_0, in_1;
  wire [67:0] z;
  CDN_bmux2 g1(.sel0 (ctl), .data0 (in_0[67]), .data1 (in_1[67]), .z
       (z[67]));
  CDN_bmux2 g2(.sel0 (ctl), .data0 (in_0[66]), .data1 (in_1[66]), .z
       (z[66]));
  CDN_bmux2 g3(.sel0 (ctl), .data0 (in_0[65]), .data1 (in_1[65]), .z
       (z[65]));
  CDN_bmux2 g4(.sel0 (ctl), .data0 (in_0[64]), .data1 (in_1[64]), .z
       (z[64]));
  CDN_bmux2 g5(.sel0 (ctl), .data0 (in_0[63]), .data1 (in_1[63]), .z
       (z[63]));
  CDN_bmux2 g6(.sel0 (ctl), .data0 (in_0[62]), .data1 (in_1[62]), .z
       (z[62]));
  CDN_bmux2 g7(.sel0 (ctl), .data0 (in_0[61]), .data1 (in_1[61]), .z
       (z[61]));
  CDN_bmux2 g8(.sel0 (ctl), .data0 (in_0[60]), .data1 (in_1[60]), .z
       (z[60]));
  CDN_bmux2 g9(.sel0 (ctl), .data0 (in_0[59]), .data1 (in_1[59]), .z
       (z[59]));
  CDN_bmux2 g10(.sel0 (ctl), .data0 (in_0[58]), .data1 (in_1[58]), .z
       (z[58]));
  CDN_bmux2 g11(.sel0 (ctl), .data0 (in_0[57]), .data1 (in_1[57]), .z
       (z[57]));
  CDN_bmux2 g12(.sel0 (ctl), .data0 (in_0[56]), .data1 (in_1[56]), .z
       (z[56]));
  CDN_bmux2 g13(.sel0 (ctl), .data0 (in_0[55]), .data1 (in_1[55]), .z
       (z[55]));
  CDN_bmux2 g14(.sel0 (ctl), .data0 (in_0[54]), .data1 (in_1[54]), .z
       (z[54]));
  CDN_bmux2 g15(.sel0 (ctl), .data0 (in_0[53]), .data1 (in_1[53]), .z
       (z[53]));
  CDN_bmux2 g16(.sel0 (ctl), .data0 (in_0[52]), .data1 (in_1[52]), .z
       (z[52]));
  CDN_bmux2 g17(.sel0 (ctl), .data0 (in_0[51]), .data1 (in_1[51]), .z
       (z[51]));
  CDN_bmux2 g18(.sel0 (ctl), .data0 (in_0[50]), .data1 (in_1[50]), .z
       (z[50]));
  CDN_bmux2 g19(.sel0 (ctl), .data0 (in_0[49]), .data1 (in_1[49]), .z
       (z[49]));
  CDN_bmux2 g20(.sel0 (ctl), .data0 (in_0[48]), .data1 (in_1[48]), .z
       (z[48]));
  CDN_bmux2 g21(.sel0 (ctl), .data0 (in_0[47]), .data1 (in_1[47]), .z
       (z[47]));
  CDN_bmux2 g22(.sel0 (ctl), .data0 (in_0[46]), .data1 (in_1[46]), .z
       (z[46]));
  CDN_bmux2 g23(.sel0 (ctl), .data0 (in_0[45]), .data1 (in_1[45]), .z
       (z[45]));
  CDN_bmux2 g24(.sel0 (ctl), .data0 (in_0[44]), .data1 (in_1[44]), .z
       (z[44]));
  CDN_bmux2 g25(.sel0 (ctl), .data0 (in_0[43]), .data1 (in_1[43]), .z
       (z[43]));
  CDN_bmux2 g26(.sel0 (ctl), .data0 (in_0[42]), .data1 (in_1[42]), .z
       (z[42]));
  CDN_bmux2 g27(.sel0 (ctl), .data0 (in_0[41]), .data1 (in_1[41]), .z
       (z[41]));
  CDN_bmux2 g28(.sel0 (ctl), .data0 (in_0[40]), .data1 (in_1[40]), .z
       (z[40]));
  CDN_bmux2 g29(.sel0 (ctl), .data0 (in_0[39]), .data1 (in_1[39]), .z
       (z[39]));
  CDN_bmux2 g30(.sel0 (ctl), .data0 (in_0[38]), .data1 (in_1[38]), .z
       (z[38]));
  CDN_bmux2 g31(.sel0 (ctl), .data0 (in_0[37]), .data1 (in_1[37]), .z
       (z[37]));
  CDN_bmux2 g32(.sel0 (ctl), .data0 (in_0[36]), .data1 (in_1[36]), .z
       (z[36]));
  CDN_bmux2 g33(.sel0 (ctl), .data0 (in_0[35]), .data1 (in_1[35]), .z
       (z[35]));
  CDN_bmux2 g34(.sel0 (ctl), .data0 (in_0[34]), .data1 (in_1[34]), .z
       (z[34]));
  CDN_bmux2 g35(.sel0 (ctl), .data0 (in_0[33]), .data1 (in_1[33]), .z
       (z[33]));
  CDN_bmux2 g36(.sel0 (ctl), .data0 (in_0[32]), .data1 (in_1[32]), .z
       (z[32]));
  CDN_bmux2 g37(.sel0 (ctl), .data0 (in_0[31]), .data1 (in_1[31]), .z
       (z[31]));
  CDN_bmux2 g38(.sel0 (ctl), .data0 (in_0[30]), .data1 (in_1[30]), .z
       (z[30]));
  CDN_bmux2 g39(.sel0 (ctl), .data0 (in_0[29]), .data1 (in_1[29]), .z
       (z[29]));
  CDN_bmux2 g40(.sel0 (ctl), .data0 (in_0[28]), .data1 (in_1[28]), .z
       (z[28]));
  CDN_bmux2 g41(.sel0 (ctl), .data0 (in_0[27]), .data1 (in_1[27]), .z
       (z[27]));
  CDN_bmux2 g42(.sel0 (ctl), .data0 (in_0[26]), .data1 (in_1[26]), .z
       (z[26]));
  CDN_bmux2 g43(.sel0 (ctl), .data0 (in_0[25]), .data1 (in_1[25]), .z
       (z[25]));
  CDN_bmux2 g44(.sel0 (ctl), .data0 (in_0[24]), .data1 (in_1[24]), .z
       (z[24]));
  CDN_bmux2 g45(.sel0 (ctl), .data0 (in_0[23]), .data1 (in_1[23]), .z
       (z[23]));
  CDN_bmux2 g46(.sel0 (ctl), .data0 (in_0[22]), .data1 (in_1[22]), .z
       (z[22]));
  CDN_bmux2 g47(.sel0 (ctl), .data0 (in_0[21]), .data1 (in_1[21]), .z
       (z[21]));
  CDN_bmux2 g48(.sel0 (ctl), .data0 (in_0[20]), .data1 (in_1[20]), .z
       (z[20]));
  CDN_bmux2 g49(.sel0 (ctl), .data0 (in_0[19]), .data1 (in_1[19]), .z
       (z[19]));
  CDN_bmux2 g50(.sel0 (ctl), .data0 (in_0[18]), .data1 (in_1[18]), .z
       (z[18]));
  CDN_bmux2 g51(.sel0 (ctl), .data0 (in_0[17]), .data1 (in_1[17]), .z
       (z[17]));
  CDN_bmux2 g52(.sel0 (ctl), .data0 (in_0[16]), .data1 (in_1[16]), .z
       (z[16]));
  CDN_bmux2 g53(.sel0 (ctl), .data0 (in_0[15]), .data1 (in_1[15]), .z
       (z[15]));
  CDN_bmux2 g54(.sel0 (ctl), .data0 (in_0[14]), .data1 (in_1[14]), .z
       (z[14]));
  CDN_bmux2 g55(.sel0 (ctl), .data0 (in_0[13]), .data1 (in_1[13]), .z
       (z[13]));
  CDN_bmux2 g56(.sel0 (ctl), .data0 (in_0[12]), .data1 (in_1[12]), .z
       (z[12]));
  CDN_bmux2 g57(.sel0 (ctl), .data0 (in_0[11]), .data1 (in_1[11]), .z
       (z[11]));
  CDN_bmux2 g58(.sel0 (ctl), .data0 (in_0[10]), .data1 (in_1[10]), .z
       (z[10]));
  CDN_bmux2 g59(.sel0 (ctl), .data0 (in_0[9]), .data1 (in_1[9]), .z
       (z[9]));
  CDN_bmux2 g60(.sel0 (ctl), .data0 (in_0[8]), .data1 (in_1[8]), .z
       (z[8]));
  CDN_bmux2 g61(.sel0 (ctl), .data0 (in_0[7]), .data1 (in_1[7]), .z
       (z[7]));
  CDN_bmux2 g62(.sel0 (ctl), .data0 (in_0[6]), .data1 (in_1[6]), .z
       (z[6]));
  CDN_bmux2 g63(.sel0 (ctl), .data0 (in_0[5]), .data1 (in_1[5]), .z
       (z[5]));
  CDN_bmux2 g64(.sel0 (ctl), .data0 (in_0[4]), .data1 (in_1[4]), .z
       (z[4]));
  CDN_bmux2 g65(.sel0 (ctl), .data0 (in_0[3]), .data1 (in_1[3]), .z
       (z[3]));
  CDN_bmux2 g66(.sel0 (ctl), .data0 (in_0[2]), .data1 (in_1[2]), .z
       (z[2]));
  CDN_bmux2 g67(.sel0 (ctl), .data0 (in_0[1]), .data1 (in_1[1]), .z
       (z[1]));
  CDN_bmux2 g68(.sel0 (ctl), .data0 (in_0[0]), .data1 (in_1[0]), .z
       (z[0]));
endmodule

module fx68k(clk, extReset, pwrUp, enPhi1, enPhi2, eRWn, ASn, LDSn,
     UDSn, E, VMAn, FC0, FC1, FC2, BGn, oRESETn, oHALTEDn, DTACKn,
     VPAn, BERRn, BRn, BGACKn, IPL0n, IPL1n, IPL2n, iEdb, oEdb, eab);
  input clk, extReset, pwrUp, enPhi1, enPhi2, DTACKn, VPAn, BERRn, BRn,
       BGACKn, IPL0n, IPL1n, IPL2n;
  input [15:0] iEdb;
  output eRWn, ASn, LDSn, UDSn, E, VMAn, FC0, FC1, FC2, BGn, oRESETn,
       oHALTEDn;
  output [15:0] oEdb;
  output [23:1] eab;
  wire clk, extReset, pwrUp, enPhi1, enPhi2, DTACKn, VPAn, BERRn, BRn,
       BGACKn, IPL0n, IPL1n, IPL2n;
  wire [15:0] iEdb;
  wire eRWn, ASn, LDSn, UDSn, E, VMAn, FC0, FC1, FC2, BGn, oRESETn,
       oHALTEDn;
  wire [15:0] oEdb;
  wire [23:1] eab;
  wire [9:0] nma;
  wire [8:0] orgAddr;
  wire [8:0] nanoAddr;
  wire [67:0] nanoOutput;
  wire [9:0] microAddr;
  wire [16:0] microOutput;
  wire [15:0] Ir;
  wire [9:0] a1;
  wire [9:0] a2;
  wire [9:0] a3;
  wire [16:0] microLatch;
  wire [2:0] pswI;
  wire [7:0] ccr;
  wire [15:0] Irc;
  wire [15:0] alue;
  wire [15:0] Ird;
  wire [3:0] tvn;
  wire [1:0] \Nanod[aluDctrl] ;
  wire [2:0] \Nanod[aluColumn] ;
  wire [1:0] \Nanod[dobCtrl] ;
  wire [2:0] \Nanod[auCntrl] ;
  wire [5:0] \Irdecod[macroTvn] ;
  wire [15:0] \Irdecod[ftuConst] ;
  wire [2:0] \Irdecod[ry] ;
  wire [2:0] \Irdecod[rx] ;
  wire [15:0] ftu;
  wire [15:0] Abl;
  wire [67:0] nanoLatch;
  wire [31:0] tState;
  wire [2:0] iIpl;
  wire [3:0] eCntr;
  wire [3:0] tvnLatch;
  wire [15:0] tvnMux;
  wire [4:0] ssw;
  wire [2:0] inl;
  wire [2:0] rIpl;
  wire A0Err, Avia, BRi, BeDebounced, BeI, BeiDelay, BerrA, BgackI;
  wire Err6591, Iac, \Irdecod[implicitSp] , \Irdecod[inhibitCcr] ,
       \Irdecod[isByte] , \Irdecod[isMovep] , \Irdecod[isPcRel] ,
       \Irdecod[isTas] ;
  wire \Irdecod[movemPreDecr] , \Irdecod[rxIsAreg] , \Irdecod[rxIsDt] ,
       \Irdecod[rxIsMovem] , \Irdecod[rxIsUsp] , \Irdecod[ryIsAreg] ,
       \Irdecod[ryIsDt] , \Irdecod[toCcr] ;
  wire \Nanod[Ir2Ird] , \Nanod[ab2Aob] , \Nanod[abd2Alub] ,
       \Nanod[abd2Dcr] , \Nanod[abdIsByte] , \Nanod[abh2Ath] ,
       \Nanod[abh2reg] , \Nanod[abh2rxh] ;
  wire \Nanod[abh2ryh] , \Nanod[abl2Atl] , \Nanod[abl2Pren] ,
       \Nanod[abl2reg] , \Nanod[abl2rxl] , \Nanod[abl2ryl] ,
       \Nanod[ablAbd] , \Nanod[ablAbh] ;
  wire \Nanod[alu2Abd] , \Nanod[alu2Dbd] , \Nanod[aluActrl] ,
       \Nanod[aluFinish] , \Nanod[aluInit] , \Nanod[alue2Dbd] ,
       \Nanod[aob2Ab] , \Nanod[ath2Abh] ;
  wire \Nanod[ath2Dbh] , \Nanod[atl2Abl] , \Nanod[atl2Dbl] ,
       \Nanod[au2Ab] , \Nanod[au2Aob] , \Nanod[au2Db] , \Nanod[au2Pc] ,
       \Nanod[auClkEn] ;
  wire \Nanod[busByte] , \Nanod[clrTpend] , \Nanod[const2Ftu] ,
       \Nanod[db2Aob] , \Nanod[dbd2Alub] , \Nanod[dbd2Alue] ,
       \Nanod[dbh2Ath] , \Nanod[dbh2reg] ;
  wire \Nanod[dbh2rxh] , \Nanod[dbh2ryh] , \Nanod[dbin2Abd] ,
       \Nanod[dbin2Dbd] , \Nanod[dbl2Atl] , \Nanod[dbl2reg] ,
       \Nanod[dbl2rxl] , \Nanod[dbl2ryl] ;
  wire \Nanod[dblDbd] , \Nanod[dblDbh] , \Nanod[dcr2Dbd] ,
       \Nanod[extAbh] , \Nanod[extDbh] , \Nanod[ftu2Abl] ,
       \Nanod[ftu2Ccr] , \Nanod[ftu2Dbl] ;
  wire \Nanod[ftu2Sr] , \Nanod[initST] , \Nanod[inl2psw] ,
       \Nanod[ird2Ftu] , \Nanod[isRmc] , \Nanod[isWrite] ,
       \Nanod[noHighByte] , \Nanod[noLowByte] ;
  wire \Nanod[noSpAlign] , \Nanod[pchabh] , \Nanod[pchdbh] ,
       \Nanod[pclabl] , \Nanod[pcldbl] , \Nanod[permStart] ,
       \Nanod[pswIToFtu] , \Nanod[reg2abh] ;
  wire \Nanod[reg2abl] , \Nanod[reg2dbh] , \Nanod[reg2dbl] ,
       \Nanod[rxh2abh] , \Nanod[rxh2dbh] , \Nanod[rxl2ab] ,
       \Nanod[rxl2db] , \Nanod[rxlDbl] ;
  wire \Nanod[ryh2abh] , \Nanod[ryh2dbh] , \Nanod[ryl2ab] ,
       \Nanod[ryl2db] , \Nanod[rz] , \Nanod[sr2Ftu] , \Nanod[ssp] ,
       \Nanod[ssw2Ftu] ;
  wire \Nanod[toIrc] , \Nanod[todbin] , \Nanod[tvn2Ftu] ,
       \Nanod[updPren] , \Nanod[updSsw] , \Nanod[updTpend] ,
       \Nanod[waitBusFinish] , Spuria;
  wire Tpend, UNCONNECTED500, UNCONNECTED501, UNCONNECTED502,
       UNCONNECTED503, UNCONNECTED504, UNCONNECTED505, UNCONNECTED506;
  wire UNCONNECTED507, UNCONNECTED508, UNCONNECTED509, UNCONNECTED510,
       UNCONNECTED511, UNCONNECTED512, UNCONNECTED513, UNCONNECTED514;
  wire UNCONNECTED515, UNCONNECTED516, UNCONNECTED517, UNCONNECTED518,
       UNCONNECTED519, UNCONNECTED520, UNCONNECTED521, UNCONNECTED522;
  wire UNCONNECTED523, UNCONNECTED524, UNCONNECTED525, UNCONNECTED526,
       UNCONNECTED527, UNCONNECTED528, UNCONNECTED529, UNCONNECTED530;
  wire UNCONNECTED531, UNCONNECTED532, UNCONNECTED533, UNCONNECTED534,
       UNCONNECTED535, UNCONNECTED536, UNCONNECTED537, UNCONNECTED538;
  wire UNCONNECTED539, UNCONNECTED540, UNCONNECTED541, UNCONNECTED542,
       UNCONNECTED543, UNCONNECTED544, UNCONNECTED545, UNCONNECTED546;
  wire UNCONNECTED547, UNCONNECTED548, UNCONNECTED549, UNCONNECTED550,
       UNCONNECTED551, UNCONNECTED552, UNCONNECTED553, UNCONNECTED554;
  wire UNCONNECTED555, UNCONNECTED556, UNCONNECTED557, UNCONNECTED558,
       UNCONNECTED559, UNCONNECTED560, UNCONNECTED561, UNCONNECTED562;
  wire UNCONNECTED563, UNCONNECTED564, UNCONNECTED565, UNCONNECTED566,
       UNCONNECTED567, UNCONNECTED568, UNCONNECTED569, UNCONNECTED570;
  wire UNCONNECTED571, UNCONNECTED572, UNCONNECTED573, UNCONNECTED574,
       UNCONNECTED575, UNCONNECTED576, UNCONNECTED577, UNCONNECTED578;
  wire UNCONNECTED579, UNCONNECTED580, UNCONNECTED581, UNCONNECTED582,
       UNCONNECTED583, UNCONNECTED584, UNCONNECTED585, UNCONNECTED586;
  wire UNCONNECTED587, UNCONNECTED588, UNCONNECTED589, UNCONNECTED590,
       UNCONNECTED591, UNCONNECTED592, UNCONNECTED593, UNCONNECTED594;
  wire UNCONNECTED595, UNCONNECTED596, UNCONNECTED597, UNCONNECTED598,
       UNCONNECTED599, UNCONNECTED600, UNCONNECTED601, UNCONNECTED602;
  wire UNCONNECTED603, UNCONNECTED604, UNCONNECTED605, UNCONNECTED606,
       UNCONNECTED607, UNCONNECTED608, UNCONNECTED609, UNCONNECTED610;
  wire UNCONNECTED611, UNCONNECTED612, UNCONNECTED613, UNCONNECTED614,
       UNCONNECTED615, UNCONNECTED616, UNCONNECTED617, UNCONNECTED618;
  wire UNCONNECTED619, UNCONNECTED620, UNCONNECTED621, UNCONNECTED622,
       UNCONNECTED623, UNCONNECTED624, UNCONNECTED625, UNCONNECTED626;
  wire UNCONNECTED627, UNCONNECTED628, UNCONNECTED629, UNCONNECTED630,
       UNCONNECTED631, UNCONNECTED632, UNCONNECTED633, UNCONNECTED634;
  wire UNCONNECTED635, UNCONNECTED636, UNCONNECTED637, UNCONNECTED638,
       UNCONNECTED639, UNCONNECTED640, UNCONNECTED641, UNCONNECTED642;
  wire UNCONNECTED643, UNCONNECTED644, UNCONNECTED645, UNCONNECTED646,
       UNCONNECTED647, UNCONNECTED648, UNCONNECTED649, UNCONNECTED650;
  wire UNCONNECTED651, UNCONNECTED652, UNCONNECTED653, UNCONNECTED654,
       UNCONNECTED655, UNCONNECTED656, UNCONNECTED657, UNCONNECTED658;
  wire UNCONNECTED659, UNCONNECTED660, UNCONNECTED661, UNCONNECTED662,
       UNCONNECTED663, UNCONNECTED664, UNCONNECTED665, UNCONNECTED666;
  wire Vpai, addrOe, aob0, au05z, bciWrite, bgBlock, busAddrErr,
       busAvail;
  wire busIsByte, busStarting, dcr4, enErrClk, enT1, enT2, enT3, enT4;
  wire excRst, iAddrErr, iBusErr, iStop, inExcept01, intPend, iplComp,
       iplStable;
  wire irdToCcr_t4, isIllegal, isLineA, isLineF, isPriv, n_601, n_602,
       n_603;
  wire n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620;
  wire n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_649, n_650;
  wire n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682;
  wire n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755;
  wire n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_783, n_784, n_801, n_802, n_803;
  wire n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811;
  wire n_813, n_815, n_817, n_818, n_822, n_824, n_825, n_827;
  wire n_828, n_830, n_831, n_833, n_843, n_844, n_845, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_866;
  wire n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874;
  wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_885;
  wire n_886, n_892, n_893, n_894, n_895, n_896, n_897, n_898;
  wire n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907;
  wire n_908, n_911, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
  wire n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934;
  wire n_935, n_936, n_937, n_938, n_939, n_940, n_945, n_946;
  wire n_947, n_948, n_954, n_955, n_956, n_957, n_1005, n_1006;
  wire n_1007, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031;
  wire n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1041, n_1042;
  wire n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050;
  wire n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058;
  wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1072, n_1073, n_1074, n_1075, n_1076, n_1654, n_1663, n_1669;
  wire n_1774, n_1777, n_1778, n_1779, n_1780, n_1781, n_1798, n_1804;
  wire n_1810, n_1811, n_1812, n_1815, n_1820, n_1825, n_1826, n_1829;
  wire n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837;
  wire n_1838, nmi, oHalted, oReset, prenEmpty, prevNmi, pswS, pswT;
  wire rAddrErr, rBerr, rDtack, rstUrom, updIll, wClk, waitBusCycle,
       xVma;
  wire ze;
  fx68k_microToNanoAddr microToNanoAddr(.uAddr (nma), .orgAddr
       (orgAddr));
  nanoRom nanoRom(.clk (clk), .nanoAddr (nanoAddr), .nanoOutput
       (nanoOutput));
  uRom uRom(.clk (clk), .microAddr (microAddr), .microOutput
       (microOutput));
  fx68k_uaddrDecode uaddrDecode(.opcode (Ir), .a1 (a1), .a2 (a2), .a3
       (a3), .isPriv (isPriv), .isIllegal (isIllegal), .isLineA
       (isLineA), .isLineF (isLineF), .lineBmap ({UNCONNECTED515,
       UNCONNECTED514, UNCONNECTED513, UNCONNECTED512, UNCONNECTED511,
       UNCONNECTED510, UNCONNECTED509, UNCONNECTED508, UNCONNECTED507,
       UNCONNECTED506, UNCONNECTED505, UNCONNECTED504, UNCONNECTED503,
       UNCONNECTED502, UNCONNECTED501, UNCONNECTED500}));
  fx68k_sequencer sequencer(.\Clks[enPhi2]  (enPhi2), .\Clks[enPhi1] 
       (enPhi1), .\Clks[pwrUp]  (pwrUp), .\Clks[extReset]  (extReset),
       .\Clks[clk]  (clk), .enT3 (enT3), .microLatch (microLatch),
       .A0Err (A0Err), .BerrA (BerrA), .busAddrErr (busAddrErr),
       .Spuria (Spuria), .Avia (Avia), .Tpend (Tpend), .intPend
       (intPend), .isIllegal (isIllegal), .isPriv (isPriv), .excRst
       (excRst), .isLineA (isLineA), .isLineF (isLineF), .psw ({pswT,
       1'b0, pswS, 2'b00, pswI, ccr}), .prenEmpty (prenEmpty), .au05z
       (au05z), .dcr4 (dcr4), .ze (ze), .i11 (Irc[11]), .alue01
       (alue[1:0]), .Ird (Ird), .a1 (a1), .a2 (a2), .a3 (a3), .tvn
       (tvn), .nma (nma));
  fx68k_excUnit excUnit(.\Clks[enPhi2]  (enPhi2), .\Clks[enPhi1] 
       (enPhi1), .\Clks[pwrUp]  (pwrUp), .\Clks[extReset]  (extReset),
       .\Clks[clk]  (clk), .enT1 (enT1), .enT2 (enT2), .enT3 (enT3),
       .enT4 (enT4), .\Nanod[abdIsByte]  (\Nanod[abdIsByte] ),
       .\Nanod[dblDbh]  (\Nanod[dblDbh] ), .\Nanod[dblDbd] 
       (\Nanod[dblDbd] ), .\Nanod[ablAbh]  (\Nanod[ablAbh] ),
       .\Nanod[ablAbd]  (\Nanod[ablAbd] ), .\Nanod[extAbh] 
       (\Nanod[extAbh] ), .\Nanod[extDbh]  (\Nanod[extDbh] ),
       .\Nanod[dbin2Dbd]  (\Nanod[dbin2Dbd] ), .\Nanod[dbin2Abd] 
       (\Nanod[dbin2Abd] ), .\Nanod[au2Pc]  (\Nanod[au2Pc] ),
       .\Nanod[au2Ab]  (\Nanod[au2Ab] ), .\Nanod[au2Db]  (\Nanod[au2Db]
       ), .\Nanod[alu2Abd]  (\Nanod[alu2Abd] ), .\Nanod[alu2Dbd] 
       (\Nanod[alu2Dbd] ), .\Nanod[abd2Alub]  (\Nanod[abd2Alub] ),
       .\Nanod[dbd2Alub]  (\Nanod[dbd2Alub] ), .\Nanod[alue2Dbd] 
       (\Nanod[alue2Dbd] ), .\Nanod[dbd2Alue]  (\Nanod[dbd2Alue] ),
       .\Nanod[dcr2Dbd]  (\Nanod[dcr2Dbd] ), .\Nanod[abd2Dcr] 
       (\Nanod[abd2Dcr] ), .\Nanod[aluFinish]  (\Nanod[aluFinish] ),
       .\Nanod[aluInit]  (\Nanod[aluInit] ), .\Nanod[aluActrl] 
       (\Nanod[aluActrl] ), .\Nanod[aluDctrl]  ({\Nanod[aluDctrl] [1],
       \Nanod[aluDctrl] [0]}), .\Nanod[aluColumn] 
       ({\Nanod[aluColumn] [2], \Nanod[aluColumn] [1],
       \Nanod[aluColumn] [0]}), .\Nanod[rxlDbl]  (\Nanod[rxlDbl] ),
       .\Nanod[rz]  (\Nanod[rz] ), .\Nanod[abl2ryl]  (\Nanod[abl2ryl]
       ), .\Nanod[dbl2ryl]  (\Nanod[dbl2ryl] ), .\Nanod[ryh2abh] 
       (\Nanod[ryh2abh] ), .\Nanod[ryh2dbh]  (\Nanod[ryh2dbh] ),
       .\Nanod[ryl2ab]  (\Nanod[ryl2ab] ), .\Nanod[ryl2db] 
       (\Nanod[ryl2db] ), .\Nanod[abh2ryh]  (\Nanod[abh2ryh] ),
       .\Nanod[dbh2ryh]  (\Nanod[dbh2ryh] ), .\Nanod[abh2rxh] 
       (\Nanod[abh2rxh] ), .\Nanod[abl2rxl]  (\Nanod[abl2rxl] ),
       .\Nanod[rxl2ab]  (\Nanod[rxl2ab] ), .\Nanod[rxl2db] 
       (\Nanod[rxl2db] ), .\Nanod[dbh2rxh]  (\Nanod[dbh2rxh] ),
       .\Nanod[dbl2rxl]  (\Nanod[dbl2rxl] ), .\Nanod[rxh2abh] 
       (\Nanod[rxh2abh] ), .\Nanod[rxh2dbh]  (\Nanod[rxh2dbh] ),
       .\Nanod[pchabh]  (\Nanod[pchabh] ), .\Nanod[pclabl] 
       (\Nanod[pclabl] ), .\Nanod[pcldbl]  (\Nanod[pcldbl] ),
       .\Nanod[pchdbh]  (\Nanod[pchdbh] ), .\Nanod[ssp]  (\Nanod[ssp]
       ), .\Nanod[reg2dbh]  (\Nanod[reg2dbh] ), .\Nanod[reg2dbl] 
       (\Nanod[reg2dbl] ), .\Nanod[dbl2reg]  (\Nanod[dbl2reg] ),
       .\Nanod[dbh2reg]  (\Nanod[dbh2reg] ), .\Nanod[reg2abh] 
       (\Nanod[reg2abh] ), .\Nanod[reg2abl]  (\Nanod[reg2abl] ),
       .\Nanod[abl2reg]  (\Nanod[abl2reg] ), .\Nanod[abh2reg] 
       (\Nanod[abh2reg] ), .\Nanod[dobCtrl]  ({\Nanod[dobCtrl] [1],
       \Nanod[dobCtrl] [0]}), .\Nanod[updSsw]  (\Nanod[updSsw] ),
       .\Nanod[aob2Ab]  (\Nanod[aob2Ab] ), .\Nanod[au2Aob] 
       (\Nanod[au2Aob] ), .\Nanod[ab2Aob]  (\Nanod[ab2Aob] ),
       .\Nanod[db2Aob]  (\Nanod[db2Aob] ), .\Nanod[ath2Abh] 
       (\Nanod[ath2Abh] ), .\Nanod[ath2Dbh]  (\Nanod[ath2Dbh] ),
       .\Nanod[dbh2Ath]  (\Nanod[dbh2Ath] ), .\Nanod[abh2Ath] 
       (\Nanod[abh2Ath] ), .\Nanod[atl2Dbl]  (\Nanod[atl2Dbl] ),
       .\Nanod[atl2Abl]  (\Nanod[atl2Abl] ), .\Nanod[abl2Atl] 
       (\Nanod[abl2Atl] ), .\Nanod[dbl2Atl]  (\Nanod[dbl2Atl] ),
       .\Nanod[toIrc]  (\Nanod[toIrc] ), .\Nanod[todbin] 
       (\Nanod[todbin] ), .\Nanod[auCntrl]  ({\Nanod[auCntrl] [2],
       \Nanod[auCntrl] [1], \Nanod[auCntrl] [0]}), .\Nanod[noSpAlign] 
       (\Nanod[noSpAlign] ), .\Nanod[auClkEn]  (\Nanod[auClkEn] ),
       .\Nanod[Ir2Ird]  (\Nanod[Ir2Ird] ), .\Nanod[initST] 
       (\Nanod[initST] ), .\Nanod[ssw2Ftu]  (\Nanod[ssw2Ftu] ),
       .\Nanod[ird2Ftu]  (\Nanod[ird2Ftu] ), .\Nanod[pswIToFtu] 
       (\Nanod[pswIToFtu] ), .\Nanod[ftu2Ccr]  (\Nanod[ftu2Ccr] ),
       .\Nanod[sr2Ftu]  (\Nanod[sr2Ftu] ), .\Nanod[ftu2Sr] 
       (\Nanod[ftu2Sr] ), .\Nanod[inl2psw]  (\Nanod[inl2psw] ),
       .\Nanod[updPren]  (\Nanod[updPren] ), .\Nanod[abl2Pren] 
       (\Nanod[abl2Pren] ), .\Nanod[ftu2Abl]  (\Nanod[ftu2Abl] ),
       .\Nanod[ftu2Dbl]  (\Nanod[ftu2Dbl] ), .\Nanod[const2Ftu] 
       (\Nanod[const2Ftu] ), .\Nanod[tvn2Ftu]  (\Nanod[tvn2Ftu] ),
       .\Nanod[clrTpend]  (\Nanod[clrTpend] ), .\Nanod[updTpend] 
       (\Nanod[updTpend] ), .\Nanod[noHighByte]  (\Nanod[noHighByte] ),
       .\Nanod[noLowByte]  (\Nanod[noLowByte] ), .\Nanod[isRmc] 
       (\Nanod[isRmc] ), .\Nanod[busByte]  (\Nanod[busByte] ),
       .\Nanod[isWrite]  (\Nanod[isWrite] ), .\Nanod[waitBusFinish] 
       (\Nanod[waitBusFinish] ), .\Nanod[permStart]  (\Nanod[permStart]
       ), .\Irdecod[inhibitCcr]  (\Irdecod[inhibitCcr] ),
       .\Irdecod[macroTvn]  ({\Irdecod[macroTvn] [5],
       \Irdecod[macroTvn] [4], \Irdecod[macroTvn] [3],
       \Irdecod[macroTvn] [2], \Irdecod[macroTvn] [1],
       \Irdecod[macroTvn] [0]}), .\Irdecod[ftuConst] 
       ({\Irdecod[ftuConst] [15], \Irdecod[ftuConst] [14],
       \Irdecod[ftuConst] [13], \Irdecod[ftuConst] [12],
       \Irdecod[ftuConst] [11], \Irdecod[ftuConst] [10],
       \Irdecod[ftuConst] [9], \Irdecod[ftuConst] [8],
       \Irdecod[ftuConst] [7], \Irdecod[ftuConst] [6],
       \Irdecod[ftuConst] [5], \Irdecod[ftuConst] [4],
       \Irdecod[ftuConst] [3], \Irdecod[ftuConst] [2],
       \Irdecod[ftuConst] [1], \Irdecod[ftuConst] [0]}),
       .\Irdecod[ryIsAreg]  (\Irdecod[ryIsAreg] ), .\Irdecod[rxIsAreg] 
       (\Irdecod[rxIsAreg] ), .\Irdecod[ry]  ({\Irdecod[ry] [2],
       \Irdecod[ry] [1], \Irdecod[ry] [0]}), .\Irdecod[rx] 
       ({\Irdecod[rx] [2], \Irdecod[rx] [1], \Irdecod[rx] [0]}),
       .\Irdecod[isMovep]  (\Irdecod[isMovep] ), .\Irdecod[isByte] 
       (\Irdecod[isByte] ), .\Irdecod[movemPreDecr] 
       (\Irdecod[movemPreDecr] ), .\Irdecod[rxIsMovem] 
       (\Irdecod[rxIsMovem] ), .\Irdecod[rxIsUsp]  (\Irdecod[rxIsUsp]
       ), .\Irdecod[ryIsDt]  (\Irdecod[ryIsDt] ), .\Irdecod[rxIsDt] 
       (\Irdecod[rxIsDt] ), .\Irdecod[toCcr]  (\Irdecod[toCcr] ),
       .\Irdecod[implicitSp]  (\Irdecod[implicitSp] ), .\Irdecod[isTas]
        (\Irdecod[isTas] ), .\Irdecod[isPcRel]  (\Irdecod[isPcRel] ),
       .Ird (Ird), .pswS (pswS), .ftu (ftu), .iEdb (iEdb), .ccr (ccr),
       .alue (alue), .prenEmpty (prenEmpty), .au05z (au05z), .dcr4
       (dcr4), .ze (ze), .aob0 (aob0), .AblOut (Abl), .Irc (Irc), .oEdb
       (oEdb), .eab (eab));
  fx68k_nDecoder3 nDecoder(.\Clks[enPhi2]  (enPhi2), .\Clks[enPhi1] 
       (enPhi1), .\Clks[pwrUp]  (pwrUp), .\Clks[extReset]  (extReset),
       .\Clks[clk]  (clk), .\Irdecod[inhibitCcr]  (\Irdecod[inhibitCcr]
       ), .\Irdecod[macroTvn]  ({\Irdecod[macroTvn] [5],
       \Irdecod[macroTvn] [4], \Irdecod[macroTvn] [3],
       \Irdecod[macroTvn] [2], \Irdecod[macroTvn] [1],
       \Irdecod[macroTvn] [0]}), .\Irdecod[ftuConst] 
       ({\Irdecod[ftuConst] [15], \Irdecod[ftuConst] [14],
       \Irdecod[ftuConst] [13], \Irdecod[ftuConst] [12],
       \Irdecod[ftuConst] [11], \Irdecod[ftuConst] [10],
       \Irdecod[ftuConst] [9], \Irdecod[ftuConst] [8],
       \Irdecod[ftuConst] [7], \Irdecod[ftuConst] [6],
       \Irdecod[ftuConst] [5], \Irdecod[ftuConst] [4],
       \Irdecod[ftuConst] [3], \Irdecod[ftuConst] [2],
       \Irdecod[ftuConst] [1], \Irdecod[ftuConst] [0]}),
       .\Irdecod[ryIsAreg]  (\Irdecod[ryIsAreg] ), .\Irdecod[rxIsAreg] 
       (\Irdecod[rxIsAreg] ), .\Irdecod[ry]  ({\Irdecod[ry] [2],
       \Irdecod[ry] [1], \Irdecod[ry] [0]}), .\Irdecod[rx] 
       ({\Irdecod[rx] [2], \Irdecod[rx] [1], \Irdecod[rx] [0]}),
       .\Irdecod[isMovep]  (\Irdecod[isMovep] ), .\Irdecod[isByte] 
       (\Irdecod[isByte] ), .\Irdecod[movemPreDecr] 
       (\Irdecod[movemPreDecr] ), .\Irdecod[rxIsMovem] 
       (\Irdecod[rxIsMovem] ), .\Irdecod[rxIsUsp]  (\Irdecod[rxIsUsp]
       ), .\Irdecod[ryIsDt]  (\Irdecod[ryIsDt] ), .\Irdecod[rxIsDt] 
       (\Irdecod[rxIsDt] ), .\Irdecod[toCcr]  (\Irdecod[toCcr] ),
       .\Irdecod[implicitSp]  (\Irdecod[implicitSp] ), .\Irdecod[isTas]
        (\Irdecod[isTas] ), .\Irdecod[isPcRel]  (\Irdecod[isPcRel] ),
       .\Nanod[abdIsByte]  (\Nanod[abdIsByte] ), .\Nanod[dblDbh] 
       (\Nanod[dblDbh] ), .\Nanod[dblDbd]  (\Nanod[dblDbd] ),
       .\Nanod[ablAbh]  (\Nanod[ablAbh] ), .\Nanod[ablAbd] 
       (\Nanod[ablAbd] ), .\Nanod[extAbh]  (\Nanod[extAbh] ),
       .\Nanod[extDbh]  (\Nanod[extDbh] ), .\Nanod[dbin2Dbd] 
       (\Nanod[dbin2Dbd] ), .\Nanod[dbin2Abd]  (\Nanod[dbin2Abd] ),
       .\Nanod[au2Pc]  (\Nanod[au2Pc] ), .\Nanod[au2Ab]  (\Nanod[au2Ab]
       ), .\Nanod[au2Db]  (\Nanod[au2Db] ), .\Nanod[alu2Abd] 
       (\Nanod[alu2Abd] ), .\Nanod[alu2Dbd]  (\Nanod[alu2Dbd] ),
       .\Nanod[abd2Alub]  (\Nanod[abd2Alub] ), .\Nanod[dbd2Alub] 
       (\Nanod[dbd2Alub] ), .\Nanod[alue2Dbd]  (\Nanod[alue2Dbd] ),
       .\Nanod[dbd2Alue]  (\Nanod[dbd2Alue] ), .\Nanod[dcr2Dbd] 
       (\Nanod[dcr2Dbd] ), .\Nanod[abd2Dcr]  (\Nanod[abd2Dcr] ),
       .\Nanod[aluFinish]  (\Nanod[aluFinish] ), .\Nanod[aluInit] 
       (\Nanod[aluInit] ), .\Nanod[aluActrl]  (\Nanod[aluActrl] ),
       .\Nanod[aluDctrl]  ({\Nanod[aluDctrl] [1], \Nanod[aluDctrl]
       [0]}), .\Nanod[aluColumn]  ({\Nanod[aluColumn] [2],
       \Nanod[aluColumn] [1], \Nanod[aluColumn] [0]}), .\Nanod[rxlDbl] 
       (\Nanod[rxlDbl] ), .\Nanod[rz]  (\Nanod[rz] ), .\Nanod[abl2ryl] 
       (\Nanod[abl2ryl] ), .\Nanod[dbl2ryl]  (\Nanod[dbl2ryl] ),
       .\Nanod[ryh2abh]  (\Nanod[ryh2abh] ), .\Nanod[ryh2dbh] 
       (\Nanod[ryh2dbh] ), .\Nanod[ryl2ab]  (\Nanod[ryl2ab] ),
       .\Nanod[ryl2db]  (\Nanod[ryl2db] ), .\Nanod[abh2ryh] 
       (\Nanod[abh2ryh] ), .\Nanod[dbh2ryh]  (\Nanod[dbh2ryh] ),
       .\Nanod[abh2rxh]  (\Nanod[abh2rxh] ), .\Nanod[abl2rxl] 
       (\Nanod[abl2rxl] ), .\Nanod[rxl2ab]  (\Nanod[rxl2ab] ),
       .\Nanod[rxl2db]  (\Nanod[rxl2db] ), .\Nanod[dbh2rxh] 
       (\Nanod[dbh2rxh] ), .\Nanod[dbl2rxl]  (\Nanod[dbl2rxl] ),
       .\Nanod[rxh2abh]  (\Nanod[rxh2abh] ), .\Nanod[rxh2dbh] 
       (\Nanod[rxh2dbh] ), .\Nanod[pchabh]  (\Nanod[pchabh] ),
       .\Nanod[pclabl]  (\Nanod[pclabl] ), .\Nanod[pcldbl] 
       (\Nanod[pcldbl] ), .\Nanod[pchdbh]  (\Nanod[pchdbh] ),
       .\Nanod[ssp]  (\Nanod[ssp] ), .\Nanod[reg2dbh]  (\Nanod[reg2dbh]
       ), .\Nanod[reg2dbl]  (\Nanod[reg2dbl] ), .\Nanod[dbl2reg] 
       (\Nanod[dbl2reg] ), .\Nanod[dbh2reg]  (\Nanod[dbh2reg] ),
       .\Nanod[reg2abh]  (\Nanod[reg2abh] ), .\Nanod[reg2abl] 
       (\Nanod[reg2abl] ), .\Nanod[abl2reg]  (\Nanod[abl2reg] ),
       .\Nanod[abh2reg]  (\Nanod[abh2reg] ), .\Nanod[dobCtrl] 
       ({\Nanod[dobCtrl] [1], \Nanod[dobCtrl] [0]}), .\Nanod[updSsw] 
       (\Nanod[updSsw] ), .\Nanod[aob2Ab]  (\Nanod[aob2Ab] ),
       .\Nanod[au2Aob]  (\Nanod[au2Aob] ), .\Nanod[ab2Aob] 
       (\Nanod[ab2Aob] ), .\Nanod[db2Aob]  (\Nanod[db2Aob] ),
       .\Nanod[ath2Abh]  (\Nanod[ath2Abh] ), .\Nanod[ath2Dbh] 
       (\Nanod[ath2Dbh] ), .\Nanod[dbh2Ath]  (\Nanod[dbh2Ath] ),
       .\Nanod[abh2Ath]  (\Nanod[abh2Ath] ), .\Nanod[atl2Dbl] 
       (\Nanod[atl2Dbl] ), .\Nanod[atl2Abl]  (\Nanod[atl2Abl] ),
       .\Nanod[abl2Atl]  (\Nanod[abl2Atl] ), .\Nanod[dbl2Atl] 
       (\Nanod[dbl2Atl] ), .\Nanod[toIrc]  (\Nanod[toIrc] ),
       .\Nanod[todbin]  (\Nanod[todbin] ), .\Nanod[auCntrl] 
       ({\Nanod[auCntrl] [2], \Nanod[auCntrl] [1], \Nanod[auCntrl]
       [0]}), .\Nanod[noSpAlign]  (\Nanod[noSpAlign] ),
       .\Nanod[auClkEn]  (\Nanod[auClkEn] ), .\Nanod[Ir2Ird] 
       (\Nanod[Ir2Ird] ), .\Nanod[initST]  (\Nanod[initST] ),
       .\Nanod[ssw2Ftu]  (\Nanod[ssw2Ftu] ), .\Nanod[ird2Ftu] 
       (\Nanod[ird2Ftu] ), .\Nanod[pswIToFtu]  (\Nanod[pswIToFtu] ),
       .\Nanod[ftu2Ccr]  (\Nanod[ftu2Ccr] ), .\Nanod[sr2Ftu] 
       (\Nanod[sr2Ftu] ), .\Nanod[ftu2Sr]  (\Nanod[ftu2Sr] ),
       .\Nanod[inl2psw]  (\Nanod[inl2psw] ), .\Nanod[updPren] 
       (\Nanod[updPren] ), .\Nanod[abl2Pren]  (\Nanod[abl2Pren] ),
       .\Nanod[ftu2Abl]  (\Nanod[ftu2Abl] ), .\Nanod[ftu2Dbl] 
       (\Nanod[ftu2Dbl] ), .\Nanod[const2Ftu]  (\Nanod[const2Ftu] ),
       .\Nanod[tvn2Ftu]  (\Nanod[tvn2Ftu] ), .\Nanod[clrTpend] 
       (\Nanod[clrTpend] ), .\Nanod[updTpend]  (\Nanod[updTpend] ),
       .\Nanod[noHighByte]  (\Nanod[noHighByte] ), .\Nanod[noLowByte] 
       (\Nanod[noLowByte] ), .\Nanod[isRmc]  (\Nanod[isRmc] ),
       .\Nanod[busByte]  (\Nanod[busByte] ), .\Nanod[isWrite] 
       (\Nanod[isWrite] ), .\Nanod[waitBusFinish] 
       (\Nanod[waitBusFinish] ), .\Nanod[permStart]  (\Nanod[permStart]
       ), .enT2 (enT2), .enT4 (enT4), .microLatch (microLatch),
       .nanoLatch (nanoLatch));
  fx68k_irdDecode irdDecode(.ird (Ird), .\Irdecod[inhibitCcr] 
       (\Irdecod[inhibitCcr] ), .\Irdecod[macroTvn] 
       ({\Irdecod[macroTvn] [5], \Irdecod[macroTvn] [4],
       \Irdecod[macroTvn] [3], \Irdecod[macroTvn] [2],
       \Irdecod[macroTvn] [1], \Irdecod[macroTvn] [0]}),
       .\Irdecod[ftuConst]  ({\Irdecod[ftuConst] [15],
       \Irdecod[ftuConst] [14], \Irdecod[ftuConst] [13],
       \Irdecod[ftuConst] [12], \Irdecod[ftuConst] [11],
       \Irdecod[ftuConst] [10], \Irdecod[ftuConst] [9],
       \Irdecod[ftuConst] [8], \Irdecod[ftuConst] [7],
       \Irdecod[ftuConst] [6], \Irdecod[ftuConst] [5],
       \Irdecod[ftuConst] [4], \Irdecod[ftuConst] [3],
       \Irdecod[ftuConst] [2], \Irdecod[ftuConst] [1],
       \Irdecod[ftuConst] [0]}), .\Irdecod[ryIsAreg] 
       (\Irdecod[ryIsAreg] ), .\Irdecod[rxIsAreg]  (\Irdecod[rxIsAreg]
       ), .\Irdecod[ry]  ({\Irdecod[ry] [2], \Irdecod[ry] [1],
       \Irdecod[ry] [0]}), .\Irdecod[rx]  ({\Irdecod[rx] [2],
       \Irdecod[rx] [1], \Irdecod[rx] [0]}), .\Irdecod[isMovep] 
       (\Irdecod[isMovep] ), .\Irdecod[isByte]  (\Irdecod[isByte] ),
       .\Irdecod[movemPreDecr]  (\Irdecod[movemPreDecr] ),
       .\Irdecod[rxIsMovem]  (\Irdecod[rxIsMovem] ), .\Irdecod[rxIsUsp]
        (\Irdecod[rxIsUsp] ), .\Irdecod[ryIsDt]  (\Irdecod[ryIsDt] ),
       .\Irdecod[rxIsDt]  (\Irdecod[rxIsDt] ), .\Irdecod[toCcr] 
       (\Irdecod[toCcr] ), .\Irdecod[implicitSp]  (\Irdecod[implicitSp]
       ), .\Irdecod[isTas]  (\Irdecod[isTas] ), .\Irdecod[isPcRel] 
       (\Irdecod[isPcRel] ));
  fx68k_busControl busControl(.\Clks[enPhi2]  (enPhi2), .\Clks[enPhi1] 
       (enPhi1), .\Clks[pwrUp]  (pwrUp), .\Clks[extReset]  (extReset),
       .\Clks[clk]  (clk), .enT1 (enT1), .enT4 (enT4), .permStart
       (\Nanod[permStart] ), .permStop (\Nanod[waitBusFinish] ), .iStop
       (iStop), .aob0 (aob0), .isWrite (\Nanod[isWrite] ), .isByte
       (busIsByte), .isRmc (\Nanod[isRmc] ), .busAvail (busAvail),
       .bgBlock (bgBlock), .busAddrErr (busAddrErr), .waitBusCycle
       (waitBusCycle), .busStarting (busStarting), .addrOe (addrOe),
       .bciWrite (bciWrite), .rDtack (rDtack), .BeDebounced
       (BeDebounced), .Vpai (Vpai), .ASn (ASn), .LDSn (LDSn), .UDSn
       (UDSn), .eRWn (eRWn));
  fx68k_busArbiter busArbiter(.\Clks[enPhi2]  (enPhi2), .\Clks[enPhi1] 
       (enPhi1), .\Clks[pwrUp]  (pwrUp), .\Clks[extReset]  (extReset),
       .\Clks[clk]  (clk), .BRi (BRi), .BgackI (BgackI), .Halti (1'b1),
       .bgBlock (bgBlock), .busAvail (busAvail), .BGn (BGn));
  fx68k_not_op_1441 g11(.A ({IPL2n, IPL1n, IPL0n}), .Z ({n_828, n_827,
       n_825}));
  fx68k_equal_unsigned_3599 eq_163_36(.A (tState), .B (3'b100), .Z
       (n_801));
  fx68k_equal_unsigned_3601 eq_166_37(.A (tState), .B (1'b0), .Z
       (n_806));
  fx68k_equal_unsigned_3603 eq_166_54(.A (tState), .B (2'b11), .Z
       (n_807));
  fx68k_equal_unsigned_3601 eq_164_36(.A (tState), .B (1'b1), .Z
       (n_804));
  fx68k_equal_unsigned_3603 eq_165_36(.A (tState), .B (2'b10), .Z
       (n_805));
  fx68k_gt_unsigned gt_401_22(.A (iIpl), .B (pswI), .Z (iplComp));
  fx68k_add_unsigned_3681 add_473_20(.A (eCntr), .B (1'b1), .Z ({n_688,
       n_687, n_686, n_685}));
  fx68k_bmux_1503 mux_rAddrErr_491_19(.ctl (n_601), .in_0 (1'b0), .in_1
       (1'b1), .z (n_603));
  fx68k_bmux_1503 mux_rAddrErr_488_7(.ctl (extReset), .in_0 (n_603),
       .in_1 (1'b0), .z (UNCONNECTED516));
  fx68k_bmux_1503 mux_rBerr_200_7(.ctl (pwrUp), .in_0 (BERRn), .in_1
       (1'b0), .z (UNCONNECTED517));
  fx68k_bmux_1503 mux_BeI_200_7(.ctl (pwrUp), .in_0 (rBerr), .in_1
       (1'b0), .z (UNCONNECTED518));
  fx68k_bmux_1503 mux_irdToCcr_t4_540_7(.ctl (pwrUp), .in_0
       (\Irdecod[toCcr] ), .in_1 (1'b0), .z (UNCONNECTED519));
  fx68k_bmux_1503 mux_updIll_427_7(.ctl (extReset), .in_0
       (microLatch[0]), .in_1 (1'b0), .z (UNCONNECTED520));
  fx68k_bmux_1766 mux_inl_427_7(.ctl (extReset), .in_0 (iIpl), .in_1
       (3'b111), .z ({UNCONNECTED523, UNCONNECTED522, UNCONNECTED521}));
  fx68k_bmux mux_tvnMux_622_22(.ctl (n_609), .in_0 ({4'b0000,
       tvnLatch}), .in_1 (Ird[7:0]), .z ({n_617, n_616, n_615, n_614,
       n_613, n_612, n_611, n_610}));
  fx68k_bmux mux_tvnMux_620_22(.ctl (n_607), .in_0 ({n_617, n_616,
       n_615, n_614, n_613, n_612, n_611, n_610}), .in_1 ({5'b00011,
       pswI}), .z ({n_625, n_624, n_623, n_622, n_621, n_620, n_619,
       n_618}));
  fx68k_bmux mux_tvnMux_618_17(.ctl (n_606), .in_0 ({n_625, n_624,
       n_623, n_622, n_621, n_620, n_619, n_618}), .in_1 (8'b00011000),
       .z ({n_633, n_632, n_631, n_630, n_629, n_628, n_627, n_626}));
  fx68k_bmux mux_tvnMux_616_7(.ctl (inExcept01), .in_0 ({2'b00,
       \Irdecod[macroTvn] [5], \Irdecod[macroTvn] [4],
       \Irdecod[macroTvn] [3], \Irdecod[macroTvn] [2],
       \Irdecod[macroTvn] [1], \Irdecod[macroTvn] [0]}), .in_1 ({n_633,
       n_632, n_631, n_630, n_629, n_628, n_627, n_626}), .z
       (tvnMux[9:2]));
  fx68k_mux_778 mux_ftu_599_11(.ctl ({\Nanod[tvn2Ftu] , \Nanod[sr2Ftu]
       , \Nanod[ird2Ftu] , \Nanod[ssw2Ftu] , \Nanod[pswIToFtu] ,
       \Nanod[const2Ftu] , \Nanod[abl2Pren] , n_649}), .in_0
       ({6'b000000, tvnMux[9:2], 2'b00}), .in_1 ({pswT, 1'b0, pswS,
       2'b00, pswI, 3'b000, ccr[4:0]}), .in_2 (Ird), .in_3
       ({11'b00000000000, ssw}), .in_4 ({12'b111111111111, pswI,
       1'b0}), .in_5 ({\Irdecod[ftuConst] [15], \Irdecod[ftuConst]
       [14], \Irdecod[ftuConst] [13], \Irdecod[ftuConst] [12],
       \Irdecod[ftuConst] [11], \Irdecod[ftuConst] [10],
       \Irdecod[ftuConst] [9], \Irdecod[ftuConst] [8],
       \Irdecod[ftuConst] [7], \Irdecod[ftuConst] [6],
       \Irdecod[ftuConst] [5], \Irdecod[ftuConst] [4],
       \Irdecod[ftuConst] [3], \Irdecod[ftuConst] [2],
       \Irdecod[ftuConst] [1], \Irdecod[ftuConst] [0]}), .in_6 (Abl),
       .in_7 (ftu), .z ({n_665, n_664, n_663, n_662, n_661, n_660,
       n_659, n_658, n_657, n_656, n_655, n_654, n_653, n_652, n_651,
       n_650}));
  fx68k_bmux_1882 mux_ftu_596_7(.ctl (pwrUp), .in_0 ({n_665, n_664,
       n_663, n_662, n_661, n_660, n_659, n_658, n_657, n_656, n_655,
       n_654, n_653, n_652, n_651, n_650}), .in_1
       (16'b0000000000000000), .z ({UNCONNECTED539, UNCONNECTED538,
       UNCONNECTED537, UNCONNECTED536, UNCONNECTED535, UNCONNECTED534,
       UNCONNECTED533, UNCONNECTED532, UNCONNECTED531, UNCONNECTED530,
       UNCONNECTED529, UNCONNECTED528, UNCONNECTED527, UNCONNECTED526,
       UNCONNECTED525, UNCONNECTED524}));
  fx68k_bmux_1503 mux_pswS_559_21(.ctl (n_605), .in_0 (1'b1), .in_1
       (ftu[13]), .z (n_666));
  fx68k_bmux_1503 mux_pswS_540_7(.ctl (pwrUp), .in_0 (n_666), .in_1
       (1'b0), .z (UNCONNECTED540));
  fx68k_bmux_1766 mux_rFC_382_7(.ctl (extReset), .in_0 ({pswS, n_669,
       n_668}), .in_1 (3'b000), .z ({UNCONNECTED543, UNCONNECTED542,
       UNCONNECTED541}));
  fx68k_bmux_1503 mux_BerrA_506_20(.ctl (n_670), .in_0 (1'b0), .in_1
       (1'b1), .z (n_672));
  fx68k_bmux_1503 mux_BerrA_503_7(.ctl (extReset), .in_0 (n_672), .in_1
       (1'b0), .z (UNCONNECTED544));
  fx68k_bmux_1503 mux_iBusErr_497_7(.ctl (extReset), .in_0 (n_673),
       .in_1 (1'b0), .z (UNCONNECTED545));
  fx68k_bmux_299 mux_microAddr_246_7(.ctl (pwrUp), .in_0 (nma), .in_1
       (10'b0000000010), .z ({UNCONNECTED555, UNCONNECTED554,
       UNCONNECTED553, UNCONNECTED552, UNCONNECTED551, UNCONNECTED550,
       UNCONNECTED549, UNCONNECTED548, UNCONNECTED547,
       UNCONNECTED546}));
  fx68k_bmux_1766 mux_microLatch_259_12(.ctl (rstUrom), .in_0
       ({microOutput[16:15], microOutput[0]}), .in_1 (3'b000), .z
       ({n_676, n_675, n_674}));
  fx68k_bmux_1894 mux_microLatch_255_7(.ctl (extReset), .in_0 ({n_676,
       n_675, microOutput[14:1], n_674}), .in_1
       (17'b00000000000000000), .z ({UNCONNECTED572, UNCONNECTED571,
       UNCONNECTED570, UNCONNECTED569, UNCONNECTED568, UNCONNECTED567,
       UNCONNECTED566, UNCONNECTED565, UNCONNECTED564, UNCONNECTED563,
       UNCONNECTED562, UNCONNECTED561, UNCONNECTED560, UNCONNECTED559,
       UNCONNECTED558, UNCONNECTED557, UNCONNECTED556}));
  fx68k_bmux_1503 mux_A0Err_522_12(.ctl (enT3), .in_0 (1'b1), .in_1
       (1'b0), .z (n_678));
  fx68k_bmux_1503 mux_A0Err_520_7(.ctl (extReset), .in_0 (n_678), .in_1
       (1'b1), .z (UNCONNECTED573));
  fx68k_bmux_1503 mux_Tpend_553_8(.ctl (\Nanod[updTpend] ), .in_0
       (1'b0), .in_1 (pswT), .z (n_679));
  fx68k_bmux_1503 mux_Tpend_540_7(.ctl (pwrUp), .in_0 (n_679), .in_1
       (1'b0), .z (UNCONNECTED574));
  fx68k_bmux_1503 mux_prevNmi_404_7(.ctl (extReset), .in_0 (nmi), .in_1
       (1'b0), .z (UNCONNECTED575));
  fx68k_bmux_1503 mux_intPend_420_19(.ctl (n_680), .in_0 (1'b0), .in_1
       (1'b1), .z (n_682));
  fx68k_bmux_1503 mux_intPend_404_7(.ctl (extReset), .in_0 (n_682),
       .in_1 (1'b0), .z (UNCONNECTED576));
  fx68k_bmux_1503 mux_excRst_515_7(.ctl (extReset), .in_0 (1'b0), .in_1
       (1'b1), .z (UNCONNECTED577));
  fx68k_bmux_1855 mux_nanoAddr_246_7(.ctl (pwrUp), .in_0 (orgAddr),
       .in_1 (9'b000000010), .z ({UNCONNECTED586, UNCONNECTED585,
       UNCONNECTED584, UNCONNECTED583, UNCONNECTED582, UNCONNECTED581,
       UNCONNECTED580, UNCONNECTED579, UNCONNECTED578}));
  fx68k_bmux_1504 mux_eCntr_470_14(.ctl (n_684), .in_0 ({n_688, n_687,
       n_686, n_685}), .in_1 (4'b0000), .z ({n_692, n_691, n_690,
       n_689}));
  fx68k_bmux_1504 mux_eCntr_464_7(.ctl (enPhi2), .in_0 (4'b0000), .in_1
       ({n_692, n_691, n_690, n_689}), .z ({n_904, n_903, n_902,
       n_900}));
  fx68k_bmux_1503 mux_rVma_476_36(.ctl (n_693), .in_0 (1'b1), .in_1
       (1'b0), .z (UNCONNECTED587));
  fx68k_bmux_1503 mux_iStop_527_7(.ctl (extReset), .in_0 (n_695), .in_1
       (1'b0), .z (UNCONNECTED588));
  fx68k_bmux_1503 mux_Err6591_527_7(.ctl (extReset), .in_0 (enErrClk),
       .in_1 (1'b0), .z (UNCONNECTED589));
  fx68k_bmux_1503 mux_179_34(.ctl (wClk), .in_0 (1'b1), .in_1 (1'b0),
       .z (n_701));
  fx68k_mux_3649 mux_tState_174_9(.ctl ({n_696, n_697, n_698, n_699,
       n_700}), .in_0 (3'b100), .in_1 (3'b010), .in_2 (3'b011), .in_3
       (3'b100), .in_4 ({2'b00, n_701}), .z ({n_704, n_703, n_702}));
  fx68k_bmux_1766 mux_tState_171_7(.ctl (pwrUp), .in_0 ({n_704, n_703,
       n_702}), .in_1 (3'b000), .z ({UNCONNECTED592, UNCONNECTED591,
       UNCONNECTED590}));
  fx68k_mux_1527 mux_E_465_8(.ctl ({n_706, n_707, n_709}), .in_0
       (1'b0), .in_1 (1'b1), .in_2 (1'b0), .z (n_710));
  fx68k_bmux_1503 mux_E_464_7(.ctl (enPhi2), .in_0 (1'b0), .in_1
       (n_710), .z (n_897));
  fx68k_bmux_1503 mux_oHalted_367_7(.ctl (pwrUp), .in_0 (n_711), .in_1
       (1'b0), .z (UNCONNECTED593));
  fx68k_bmux_1503 mux_oReset_367_7(.ctl (pwrUp), .in_0 (n_712), .in_1
       (1'b0), .z (UNCONNECTED594));
  fx68k_bmux_1766 mux_pswI_559_21(.ctl (n_605), .in_0 (inl), .in_1
       (ftu[10:8]), .z ({n_715, n_714, n_713}));
  fx68k_bmux_1766 mux_pswI_540_7(.ctl (pwrUp), .in_0 ({n_715, n_714,
       n_713}), .in_1 (3'b000), .z ({UNCONNECTED597, UNCONNECTED596,
       UNCONNECTED595}));
  fx68k_bmux_1503 mux_pswT_559_21(.ctl (n_605), .in_0 (1'b0), .in_1
       (ftu[15]), .z (n_716));
  fx68k_bmux_1503 mux_pswT_540_7(.ctl (pwrUp), .in_0 (n_716), .in_1
       (1'b0), .z (UNCONNECTED598));
  fx68k_bmux_3758 mux_nanoLatch_259_12(.ctl (rstUrom), .in_0
       (nanoOutput), .in_1
       (68'b00000000000000000000000000000000000000000000000000000000000000000000),
       .z ({n_784, n_783, n_782, n_781, n_780, n_779, n_778, n_777,
       n_776, n_775, n_774, n_773, n_772, n_771, n_770, n_769, n_768,
       n_767, n_766, n_765, n_764, n_763, n_762, n_761, n_760, n_759,
       n_758, n_757, n_756, n_755, n_754, n_753, n_752, n_751, n_750,
       n_749, n_748, n_747, n_746, n_745, n_744, n_743, n_742, n_741,
       n_740, n_739, n_738, n_737, n_736, n_735, n_734, n_733, n_732,
       n_731, n_730, n_729, n_728, n_727, n_726, n_725, n_724, n_723,
       n_722, n_721, n_720, n_719, n_718, n_717}));
  fx68k_bmux_3758 mux_nanoLatch_255_7(.ctl (extReset), .in_0 ({n_784,
       n_783, n_782, n_781, n_780, n_779, n_778, n_777, n_776, n_775,
       n_774, n_773, n_772, n_771, n_770, n_769, n_768, n_767, n_766,
       n_765, n_764, n_763, n_762, n_761, n_760, n_759, n_758, n_757,
       n_756, n_755, n_754, n_753, n_752, n_751, n_750, n_749, n_748,
       n_747, n_746, n_745, n_744, n_743, n_742, n_741, n_740, n_739,
       n_738, n_737, n_736, n_735, n_734, n_733, n_732, n_731, n_730,
       n_729, n_728, n_727, n_726, n_725, n_724, n_723, n_722, n_721,
       n_720, n_719, n_718, n_717}), .in_1
       (68'b00000000000000000000000000000000000000000000000000000000000000000000),
       .z ({UNCONNECTED666, UNCONNECTED665, UNCONNECTED664,
       UNCONNECTED663, UNCONNECTED662, UNCONNECTED661, UNCONNECTED660,
       UNCONNECTED659, UNCONNECTED658, UNCONNECTED657, UNCONNECTED656,
       UNCONNECTED655, UNCONNECTED654, UNCONNECTED653, UNCONNECTED652,
       UNCONNECTED651, UNCONNECTED650, UNCONNECTED649, UNCONNECTED648,
       UNCONNECTED647, UNCONNECTED646, UNCONNECTED645, UNCONNECTED644,
       UNCONNECTED643, UNCONNECTED642, UNCONNECTED641, UNCONNECTED640,
       UNCONNECTED639, UNCONNECTED638, UNCONNECTED637, UNCONNECTED636,
       UNCONNECTED635, UNCONNECTED634, UNCONNECTED633, UNCONNECTED632,
       UNCONNECTED631, UNCONNECTED630, UNCONNECTED629, UNCONNECTED628,
       UNCONNECTED627, UNCONNECTED626, UNCONNECTED625, UNCONNECTED624,
       UNCONNECTED623, UNCONNECTED622, UNCONNECTED621, UNCONNECTED620,
       UNCONNECTED619, UNCONNECTED618, UNCONNECTED617, UNCONNECTED616,
       UNCONNECTED615, UNCONNECTED614, UNCONNECTED613, UNCONNECTED612,
       UNCONNECTED611, UNCONNECTED610, UNCONNECTED609, UNCONNECTED608,
       UNCONNECTED607, UNCONNECTED606, UNCONNECTED605, UNCONNECTED604,
       UNCONNECTED603, UNCONNECTED602, UNCONNECTED601, UNCONNECTED600,
       UNCONNECTED599}));
  and g1 (n_802, enPhi1, n_801);
  not g2 (n_803, wClk);
  and g3 (enT1, n_802, n_803);
  and g4 (enT2, enPhi2, n_804);
  and g5 (enT3, enPhi1, n_805);
  or g6 (n_808, n_806, n_807);
  and g7 (enT4, enPhi2, n_808);
  or g9 (n_818, BeI, BeiDelay);
  not g10 (BeDebounced, n_818);
  or g27 (n_853, \Irdecod[isByte] , \Irdecod[isMovep] );
  and g28 (busIsByte, \Nanod[busByte] , n_853);
  and g29 (iAddrErr, rAddrErr, addrOe);
  and g30 (rstUrom, enPhi1, enErrClk);
  and g34 (n_712, n_854, n_855);
  and g35 (n_711, n_856, n_855);
  and g38 (n_667, enT1, \Nanod[permStart] );
  not g39 (n_857, microLatch[15]);
  not g40 (n_858, \Irdecod[isPcRel] );
  and g41 (n_859, n_857, n_858);
  or g42 (n_669, microLatch[16], n_859);
  and g44 (n_861, n_860, \Irdecod[isPcRel] );
  or g45 (n_668, microLatch[15], n_861);
  not g47 (n_862, prevNmi);
  and g48 (n_863, nmi, n_862);
  or g49 (n_864, n_863, iplComp);
  and g50 (n_680, iplStable, n_864);
  and g53 (n_867, iplStable, n_866);
  and g55 (n_870, n_867, n_868);
  or g56 (n_681, n_869, n_870);
  and g57 (n_608, enT1, updIll);
  not g58 (n_871, BeiDelay);
  and g59 (n_877, n_871, Iac);
  not g60 (n_872, Vpai);
  and g61 (n_878, n_872, Iac);
  or g68 (enErrClk, iAddrErr, iBusErr);
  not g69 (n_881, BeI);
  not g73 (n_885, VMAn);
  and g74 (xVma, n_885, n_886);
  and g83 (n_601, busAddrErr, addrOe);
  not g84 (n_602, addrOe);
  and g85 (n_907, BerrA, n_881);
  and g87 (n_673, n_907, n_908);
  and g90 (n_911, n_881, n_908);
  and g91 (n_670, n_911, addrOe);
  and g92 (n_671, BeI, busStarting);
  and g93 (n_683, enT2, \Nanod[permStart] );
  or g95 (n_913, busAddrErr, BerrA);
  and g96 (n_677, rstUrom, n_913);
  not g97 (n_914, rBerr);
  or g98 (n_915, iAddrErr, n_914);
  and g99 (n_916, Vpai, n_915);
  or g100 (n_695, xVma, n_916);
  and g109 (n_605, \Nanod[ftu2Sr] , n_930);
  and g115 (n_634, \Nanod[updSsw] , enT3);
  not g116 (n_956, bciWrite);
  and g117 (n_705, enT1, \Nanod[Ir2Ird] );
  not g122 (n_822, pwrUp);
  not g123 (n_830, enPhi2);
  not g124 (n_917, enPhi1);
  not g126 (n_919, extReset);
  not g127 (n_926, n_601);
  not g129 (n_849, \Nanod[Ir2Ird] );
  not g131 (n_879, enT4);
  not g133 (n_936, n_605);
  not g143 (n_922, n_670);
  not g145 (n_843, rstUrom);
  not g147 (n_931, \Nanod[updTpend] );
  not g149 (n_873, n_680);
  not g153 (n_905, n_693);
  or g157 (n_708, n_706, n_707);
  not g158 (n_709, n_708);
  and g159 (n_810, enPhi2, n_696);
  and g160 (n_809, enPhi2, n_697);
  and g162 (n_811, enPhi1, n_698);
  and g164 (n_813, enPhi2, n_699);
  and g166 (n_815, enPhi1, n_700);
  and g168 (n_824, enPhi2, n_822);
  and g171 (n_831, enPhi1, n_830);
  and g172 (n_833, n_831, n_822);
  and g180 (n_844, enT3, n_843);
  or g181 (n_845, n_844, rstUrom);
  and g185 (n_850, microLatch[0], n_849);
  and g186 (n_851, n_850, enT1);
  and g187 (n_852, \Nanod[Ir2Ird] , enT1);
  and g188 (n_874, n_681, n_873);
  or g189 (n_875, n_874, n_680);
  and g190 (n_876, n_875, enPhi2);
  and g191 (n_880, n_608, n_879);
  or g192 (n_893, n_707, n_706);
  and g193 (n_892, pwrUp, n_709);
  or g194 (n_894, n_892, n_893);
  and g195 (n_896, n_894, enPhi2);
  and g196 (n_895, pwrUp, n_830);
  or g197 (n_898, n_895, n_896);
  or g199 (n_901, n_895, enPhi2);
  and g201 (n_918, enPhi2, n_917);
  and g202 (n_920, enT3, n_919);
  and g203 (n_921, n_683, n_919);
  and g204 (n_923, n_671, n_922);
  or g205 (n_924, n_923, n_670);
  and g206 (n_925, n_924, enPhi2);
  and g207 (n_927, n_602, n_926);
  or g208 (n_928, n_927, n_601);
  and g209 (n_929, n_928, enPhi1);
  and g210 (n_932, \Nanod[clrTpend] , n_931);
  or g211 (n_933, n_932, \Nanod[updTpend] );
  and g212 (n_934, n_933, enT3);
  and g213 (n_935, n_934, n_879);
  and g214 (n_937, \Nanod[initST] , n_936);
  or g215 (n_938, n_937, n_605);
  and g216 (n_939, n_938, enT3);
  and g217 (n_940, n_939, n_879);
  and g222 (n_945, \Nanod[inl2psw] , n_936);
  or g223 (n_946, n_945, n_605);
  and g224 (n_947, n_946, enT3);
  and g225 (n_948, n_947, n_879);
  and g232 (n_955, n_954, enT3);
  nor g240 (n_1006, \Nanod[tvn2Ftu] , \Nanod[sr2Ftu] , \Nanod[ird2Ftu]
       , \Nanod[ssw2Ftu] );
  nor g241 (n_1005, \Nanod[pswIToFtu] , \Nanod[const2Ftu] ,
       \Nanod[abl2Pren] );
  nand g242 (n_1007, n_1005, n_1006);
  not g243 (n_649, n_1007);
  not g244 (n_1009, tState[31]);
  not g245 (n_1010, tState[30]);
  not g246 (n_1011, tState[29]);
  not g247 (n_1012, tState[28]);
  not g248 (n_1013, tState[27]);
  not g249 (n_1014, tState[26]);
  not g250 (n_1015, tState[25]);
  not g251 (n_1016, tState[24]);
  not g252 (n_1017, tState[23]);
  not g253 (n_1018, tState[22]);
  not g254 (n_1019, tState[21]);
  not g255 (n_1020, tState[20]);
  not g256 (n_1021, tState[19]);
  not g257 (n_1022, tState[18]);
  not g258 (n_1023, tState[17]);
  not g259 (n_1024, tState[16]);
  not g260 (n_1025, tState[15]);
  not g261 (n_1026, tState[14]);
  not g262 (n_1027, tState[13]);
  not g263 (n_1028, tState[12]);
  not g264 (n_1029, tState[11]);
  not g265 (n_1030, tState[10]);
  not g266 (n_1031, tState[9]);
  not g267 (n_1032, tState[8]);
  not g268 (n_1033, tState[7]);
  not g269 (n_1034, tState[6]);
  not g270 (n_1035, tState[5]);
  not g271 (n_1036, tState[4]);
  not g272 (n_1037, tState[3]);
  nand g276 (n_1044, n_1009, n_1010, n_1011, n_1012);
  nand g277 (n_1045, n_1013, n_1014, n_1015, n_1016);
  nand g278 (n_1046, n_1017, n_1018, n_1019, n_1020);
  nand g279 (n_1047, n_1021, n_1022, n_1023, n_1024);
  nand g280 (n_1048, n_1025, n_1026, n_1027, n_1028);
  nand g281 (n_1049, n_1029, n_1030, n_1031, n_1032);
  nand g282 (n_1050, n_1033, n_1034, n_1035, n_1036);
  nand g283 (n_1051, n_1037, n_1041, n_1042, n_1043);
  nor g284 (n_1053, n_1044, n_1045, n_1046, n_1047);
  nor g285 (n_1052, n_1048, n_1049, n_1050, n_1051);
  nand g286 (n_1062, n_1052, n_1053);
  nand g287 (n_1054, n_1037, n_1041, n_1042, tState[0]);
  nor g288 (n_1055, n_1048, n_1049, n_1050, n_1054);
  nand g289 (n_1063, n_1055, n_1053);
  nand g290 (n_1056, n_1037, n_1041, tState[1], n_1043);
  nor g291 (n_1057, n_1048, n_1049, n_1050, n_1056);
  nand g292 (n_1064, n_1057, n_1053);
  nand g293 (n_1058, n_1037, n_1041, tState[1], tState[0]);
  nor g294 (n_1059, n_1048, n_1049, n_1050, n_1058);
  nand g295 (n_1065, n_1059, n_1053);
  nand g296 (n_1060, n_1037, tState[2], n_1042, n_1043);
  nor g297 (n_1061, n_1048, n_1049, n_1050, n_1060);
  nand g298 (n_1066, n_1061, n_1053);
  not g299 (n_696, n_1062);
  not g300 (n_697, n_1063);
  not g301 (n_698, n_1064);
  not g302 (n_699, n_1065);
  not g303 (n_700, n_1066);
  not g307 (n_1041, tState[2]);
  not g308 (n_1042, tState[1]);
  not g309 (n_1043, tState[0]);
  not g312 (n_1072, eCntr[1]);
  nand g313 (n_1075, eCntr[3], n_1073, n_1072, eCntr[0]);
  nand g314 (n_1076, n_1074, eCntr[2], n_1072, eCntr[0]);
  not g315 (n_706, n_1075);
  not g316 (n_707, n_1076);
  not g318 (n_1073, eCntr[2]);
  not g319 (n_1074, eCntr[3]);
  CDN_flop \tState_reg[0] (.clk (clk), .d (n_702), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[0]));
  CDN_flop \tState_reg[1] (.clk (clk), .d (n_703), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[1]));
  CDN_flop \tState_reg[2] (.clk (clk), .d (n_704), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[2]));
  CDN_flop \tState_reg[3] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[3]));
  CDN_flop \tState_reg[4] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[4]));
  CDN_flop \tState_reg[5] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[5]));
  CDN_flop \tState_reg[6] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[6]));
  CDN_flop \tState_reg[7] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[7]));
  CDN_flop \tState_reg[8] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[8]));
  CDN_flop \tState_reg[9] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (tState[9]));
  CDN_flop \tState_reg[10] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[10]));
  CDN_flop \tState_reg[11] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[11]));
  CDN_flop \tState_reg[12] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[12]));
  CDN_flop \tState_reg[13] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[13]));
  CDN_flop \tState_reg[14] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[14]));
  CDN_flop \tState_reg[15] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[15]));
  CDN_flop \tState_reg[16] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[16]));
  CDN_flop \tState_reg[17] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[17]));
  CDN_flop \tState_reg[18] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[18]));
  CDN_flop \tState_reg[19] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[19]));
  CDN_flop \tState_reg[20] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[20]));
  CDN_flop \tState_reg[21] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[21]));
  CDN_flop \tState_reg[22] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[22]));
  CDN_flop \tState_reg[23] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[23]));
  CDN_flop \tState_reg[24] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[24]));
  CDN_flop \tState_reg[25] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[25]));
  CDN_flop \tState_reg[26] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[26]));
  CDN_flop \tState_reg[27] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[27]));
  CDN_flop \tState_reg[28] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[28]));
  CDN_flop \tState_reg[29] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[29]));
  CDN_flop \tState_reg[30] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[30]));
  CDN_flop \tState_reg[31] (.clk (clk), .d (1'b0), .sena (n_817), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (tState[31]));
  CDN_flop rDtack_reg(.clk (clk), .d (DTACKn), .sena (n_824), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (rDtack));
  CDN_flop rBerr_reg(.clk (clk), .d (BERRn), .sena (enPhi2), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (rBerr));
  CDN_flop \rIpl_reg[0] (.clk (clk), .d (n_825), .sena (n_824), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (rIpl[0]));
  CDN_flop \rIpl_reg[1] (.clk (clk), .d (n_827), .sena (n_824), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (rIpl[1]));
  CDN_flop \rIpl_reg[2] (.clk (clk), .d (n_828), .sena (n_824), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (rIpl[2]));
  CDN_flop \iIpl_reg[0] (.clk (clk), .d (rIpl[0]), .sena (n_824), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (iIpl[0]));
  CDN_flop \iIpl_reg[1] (.clk (clk), .d (rIpl[1]), .sena (n_824), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (iIpl[1]));
  CDN_flop \iIpl_reg[2] (.clk (clk), .d (rIpl[2]), .sena (n_824), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (iIpl[2]));
  CDN_flop Vpai_reg(.clk (clk), .d (VPAn), .sena (n_833), .aclr (1'b0),
       .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Vpai));
  CDN_flop BeI_reg(.clk (clk), .d (rBerr), .sena (n_831), .aclr (1'b0),
       .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (BeI));
  CDN_flop BRi_reg(.clk (clk), .d (BRn), .sena (n_833), .aclr (1'b0),
       .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (BRi));
  CDN_flop BgackI_reg(.clk (clk), .d (BGACKn), .sena (n_833), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (BgackI));
  CDN_flop BeiDelay_reg(.clk (clk), .d (BeI), .sena (n_833), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (BeiDelay));
  CDN_flop \nanoLatch_reg[0] (.clk (clk), .d (n_717), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[0]));
  CDN_flop \nanoLatch_reg[1] (.clk (clk), .d (n_718), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[1]));
  CDN_flop \nanoLatch_reg[2] (.clk (clk), .d (n_719), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[2]));
  CDN_flop \nanoLatch_reg[3] (.clk (clk), .d (n_720), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[3]));
  CDN_flop \nanoLatch_reg[4] (.clk (clk), .d (n_721), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[4]));
  CDN_flop \nanoLatch_reg[5] (.clk (clk), .d (n_722), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[5]));
  CDN_flop \nanoLatch_reg[6] (.clk (clk), .d (n_723), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[6]));
  CDN_flop \nanoLatch_reg[7] (.clk (clk), .d (n_724), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[7]));
  CDN_flop \nanoLatch_reg[8] (.clk (clk), .d (n_725), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[8]));
  CDN_flop \nanoLatch_reg[9] (.clk (clk), .d (n_726), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[9]));
  CDN_flop \nanoLatch_reg[10] (.clk (clk), .d (n_727), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[10]));
  CDN_flop \nanoLatch_reg[11] (.clk (clk), .d (n_728), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[11]));
  CDN_flop \nanoLatch_reg[12] (.clk (clk), .d (n_729), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[12]));
  CDN_flop \nanoLatch_reg[13] (.clk (clk), .d (n_730), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[13]));
  CDN_flop \nanoLatch_reg[14] (.clk (clk), .d (n_731), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[14]));
  CDN_flop \nanoLatch_reg[15] (.clk (clk), .d (n_732), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[15]));
  CDN_flop \nanoLatch_reg[16] (.clk (clk), .d (n_733), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[16]));
  CDN_flop \nanoLatch_reg[17] (.clk (clk), .d (n_734), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[17]));
  CDN_flop \nanoLatch_reg[18] (.clk (clk), .d (n_735), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[18]));
  CDN_flop \nanoLatch_reg[19] (.clk (clk), .d (n_736), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[19]));
  CDN_flop \nanoLatch_reg[20] (.clk (clk), .d (n_737), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[20]));
  CDN_flop \nanoLatch_reg[21] (.clk (clk), .d (n_738), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[21]));
  CDN_flop \nanoLatch_reg[22] (.clk (clk), .d (n_739), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[22]));
  CDN_flop \nanoLatch_reg[23] (.clk (clk), .d (n_740), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[23]));
  CDN_flop \nanoLatch_reg[24] (.clk (clk), .d (n_741), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[24]));
  CDN_flop \nanoLatch_reg[25] (.clk (clk), .d (n_742), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[25]));
  CDN_flop \nanoLatch_reg[26] (.clk (clk), .d (n_743), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[26]));
  CDN_flop \nanoLatch_reg[27] (.clk (clk), .d (n_744), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[27]));
  CDN_flop \nanoLatch_reg[28] (.clk (clk), .d (n_745), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[28]));
  CDN_flop \nanoLatch_reg[29] (.clk (clk), .d (n_746), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[29]));
  CDN_flop \nanoLatch_reg[30] (.clk (clk), .d (n_747), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[30]));
  CDN_flop \nanoLatch_reg[31] (.clk (clk), .d (n_748), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[31]));
  CDN_flop \nanoLatch_reg[32] (.clk (clk), .d (n_749), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[32]));
  CDN_flop \nanoLatch_reg[33] (.clk (clk), .d (n_750), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[33]));
  CDN_flop \nanoLatch_reg[34] (.clk (clk), .d (n_751), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[34]));
  CDN_flop \nanoLatch_reg[35] (.clk (clk), .d (n_752), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[35]));
  CDN_flop \nanoLatch_reg[36] (.clk (clk), .d (n_753), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[36]));
  CDN_flop \nanoLatch_reg[37] (.clk (clk), .d (n_754), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[37]));
  CDN_flop \nanoLatch_reg[38] (.clk (clk), .d (n_755), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[38]));
  CDN_flop \nanoLatch_reg[39] (.clk (clk), .d (n_756), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[39]));
  CDN_flop \nanoLatch_reg[40] (.clk (clk), .d (n_757), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[40]));
  CDN_flop \nanoLatch_reg[41] (.clk (clk), .d (n_758), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[41]));
  CDN_flop \nanoLatch_reg[42] (.clk (clk), .d (n_759), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[42]));
  CDN_flop \nanoLatch_reg[43] (.clk (clk), .d (n_760), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[43]));
  CDN_flop \nanoLatch_reg[44] (.clk (clk), .d (n_761), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[44]));
  CDN_flop \nanoLatch_reg[45] (.clk (clk), .d (n_762), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[45]));
  CDN_flop \nanoLatch_reg[46] (.clk (clk), .d (n_763), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[46]));
  CDN_flop \nanoLatch_reg[47] (.clk (clk), .d (n_764), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[47]));
  CDN_flop \nanoLatch_reg[48] (.clk (clk), .d (n_765), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[48]));
  CDN_flop \nanoLatch_reg[49] (.clk (clk), .d (n_766), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[49]));
  CDN_flop \nanoLatch_reg[50] (.clk (clk), .d (n_767), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[50]));
  CDN_flop \nanoLatch_reg[51] (.clk (clk), .d (n_768), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[51]));
  CDN_flop \nanoLatch_reg[52] (.clk (clk), .d (n_769), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[52]));
  CDN_flop \nanoLatch_reg[53] (.clk (clk), .d (n_770), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[53]));
  CDN_flop \nanoLatch_reg[54] (.clk (clk), .d (n_771), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[54]));
  CDN_flop \nanoLatch_reg[55] (.clk (clk), .d (n_772), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[55]));
  CDN_flop \nanoLatch_reg[56] (.clk (clk), .d (n_773), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[56]));
  CDN_flop \nanoLatch_reg[57] (.clk (clk), .d (n_774), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[57]));
  CDN_flop \nanoLatch_reg[58] (.clk (clk), .d (n_775), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[58]));
  CDN_flop \nanoLatch_reg[59] (.clk (clk), .d (n_776), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[59]));
  CDN_flop \nanoLatch_reg[60] (.clk (clk), .d (n_777), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[60]));
  CDN_flop \nanoLatch_reg[61] (.clk (clk), .d (n_778), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[61]));
  CDN_flop \nanoLatch_reg[62] (.clk (clk), .d (n_779), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[62]));
  CDN_flop \nanoLatch_reg[63] (.clk (clk), .d (n_780), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[63]));
  CDN_flop \nanoLatch_reg[64] (.clk (clk), .d (n_781), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[64]));
  CDN_flop \nanoLatch_reg[65] (.clk (clk), .d (n_782), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[65]));
  CDN_flop \nanoLatch_reg[66] (.clk (clk), .d (n_783), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[66]));
  CDN_flop \nanoLatch_reg[67] (.clk (clk), .d (n_784), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (nanoLatch[67]));
  CDN_flop \microLatch_reg[0] (.clk (clk), .d (n_674), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (microLatch[0]));
  CDN_flop \microLatch_reg[1] (.clk (clk), .d (microOutput[1]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[1]));
  CDN_flop \microLatch_reg[2] (.clk (clk), .d (microOutput[2]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[2]));
  CDN_flop \microLatch_reg[3] (.clk (clk), .d (microOutput[3]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[3]));
  CDN_flop \microLatch_reg[4] (.clk (clk), .d (microOutput[4]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[4]));
  CDN_flop \microLatch_reg[5] (.clk (clk), .d (microOutput[5]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[5]));
  CDN_flop \microLatch_reg[6] (.clk (clk), .d (microOutput[6]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[6]));
  CDN_flop \microLatch_reg[7] (.clk (clk), .d (microOutput[7]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[7]));
  CDN_flop \microLatch_reg[8] (.clk (clk), .d (microOutput[8]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[8]));
  CDN_flop \microLatch_reg[9] (.clk (clk), .d (microOutput[9]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[9]));
  CDN_flop \microLatch_reg[10] (.clk (clk), .d (microOutput[10]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[10]));
  CDN_flop \microLatch_reg[11] (.clk (clk), .d (microOutput[11]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[11]));
  CDN_flop \microLatch_reg[12] (.clk (clk), .d (microOutput[12]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[12]));
  CDN_flop \microLatch_reg[13] (.clk (clk), .d (microOutput[13]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[13]));
  CDN_flop \microLatch_reg[14] (.clk (clk), .d (microOutput[14]), .sena
       (n_844), .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd
       (1'b0), .q (microLatch[14]));
  CDN_flop \microLatch_reg[15] (.clk (clk), .d (n_675), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (microLatch[15]));
  CDN_flop \microLatch_reg[16] (.clk (clk), .d (n_676), .sena (n_845),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (microLatch[16]));
  CDN_flop \microAddr_reg[0] (.clk (clk), .d (nma[0]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[0]));
  CDN_flop \microAddr_reg[1] (.clk (clk), .d (nma[1]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b1), .q
       (microAddr[1]));
  CDN_flop \microAddr_reg[2] (.clk (clk), .d (nma[2]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[2]));
  CDN_flop \microAddr_reg[3] (.clk (clk), .d (nma[3]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[3]));
  CDN_flop \microAddr_reg[4] (.clk (clk), .d (nma[4]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[4]));
  CDN_flop \microAddr_reg[5] (.clk (clk), .d (nma[5]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[5]));
  CDN_flop \microAddr_reg[6] (.clk (clk), .d (nma[6]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[6]));
  CDN_flop \microAddr_reg[7] (.clk (clk), .d (nma[7]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[7]));
  CDN_flop \microAddr_reg[8] (.clk (clk), .d (nma[8]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[8]));
  CDN_flop \microAddr_reg[9] (.clk (clk), .d (nma[9]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (microAddr[9]));
  CDN_flop \nanoAddr_reg[0] (.clk (clk), .d (orgAddr[0]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[0]));
  CDN_flop \nanoAddr_reg[1] (.clk (clk), .d (orgAddr[1]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b1), .q
       (nanoAddr[1]));
  CDN_flop \nanoAddr_reg[2] (.clk (clk), .d (orgAddr[2]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[2]));
  CDN_flop \nanoAddr_reg[3] (.clk (clk), .d (orgAddr[3]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[3]));
  CDN_flop \nanoAddr_reg[4] (.clk (clk), .d (orgAddr[4]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[4]));
  CDN_flop \nanoAddr_reg[5] (.clk (clk), .d (orgAddr[5]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[5]));
  CDN_flop \nanoAddr_reg[6] (.clk (clk), .d (orgAddr[6]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[6]));
  CDN_flop \nanoAddr_reg[7] (.clk (clk), .d (orgAddr[7]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[7]));
  CDN_flop \nanoAddr_reg[8] (.clk (clk), .d (orgAddr[8]), .sena (enT1),
       .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q
       (nanoAddr[8]));
  CDN_flop \Ir_reg[0] (.clk (clk), .d (Irc[0]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[0]));
  CDN_flop \Ir_reg[1] (.clk (clk), .d (Irc[1]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[1]));
  CDN_flop \Ir_reg[2] (.clk (clk), .d (Irc[2]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[2]));
  CDN_flop \Ir_reg[3] (.clk (clk), .d (Irc[3]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[3]));
  CDN_flop \Ir_reg[4] (.clk (clk), .d (Irc[4]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[4]));
  CDN_flop \Ir_reg[5] (.clk (clk), .d (Irc[5]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[5]));
  CDN_flop \Ir_reg[6] (.clk (clk), .d (Irc[6]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[6]));
  CDN_flop \Ir_reg[7] (.clk (clk), .d (Irc[7]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[7]));
  CDN_flop \Ir_reg[8] (.clk (clk), .d (Irc[8]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[8]));
  CDN_flop \Ir_reg[9] (.clk (clk), .d (Irc[9]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[9]));
  CDN_flop \Ir_reg[10] (.clk (clk), .d (Irc[10]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[10]));
  CDN_flop \Ir_reg[11] (.clk (clk), .d (Irc[11]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[11]));
  CDN_flop \Ir_reg[12] (.clk (clk), .d (Irc[12]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[12]));
  CDN_flop \Ir_reg[13] (.clk (clk), .d (Irc[13]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[13]));
  CDN_flop \Ir_reg[14] (.clk (clk), .d (Irc[14]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[14]));
  CDN_flop \Ir_reg[15] (.clk (clk), .d (Irc[15]), .sena (n_851), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ir[15]));
  CDN_flop \Ird_reg[0] (.clk (clk), .d (Ir[0]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[0]));
  CDN_flop \Ird_reg[1] (.clk (clk), .d (Ir[1]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[1]));
  CDN_flop \Ird_reg[2] (.clk (clk), .d (Ir[2]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[2]));
  CDN_flop \Ird_reg[3] (.clk (clk), .d (Ir[3]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[3]));
  CDN_flop \Ird_reg[4] (.clk (clk), .d (Ir[4]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[4]));
  CDN_flop \Ird_reg[5] (.clk (clk), .d (Ir[5]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[5]));
  CDN_flop \Ird_reg[6] (.clk (clk), .d (Ir[6]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[6]));
  CDN_flop \Ird_reg[7] (.clk (clk), .d (Ir[7]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[7]));
  CDN_flop \Ird_reg[8] (.clk (clk), .d (Ir[8]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[8]));
  CDN_flop \Ird_reg[9] (.clk (clk), .d (Ir[9]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[9]));
  CDN_flop \Ird_reg[10] (.clk (clk), .d (Ir[10]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[10]));
  CDN_flop \Ird_reg[11] (.clk (clk), .d (Ir[11]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[11]));
  CDN_flop \Ird_reg[12] (.clk (clk), .d (Ir[12]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[12]));
  CDN_flop \Ird_reg[13] (.clk (clk), .d (Ir[13]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[13]));
  CDN_flop \Ird_reg[14] (.clk (clk), .d (Ir[14]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[14]));
  CDN_flop \Ird_reg[15] (.clk (clk), .d (Ir[15]), .sena (n_852), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Ird[15]));
  not g627 (oRESETn, oReset);
  not g628 (oHALTEDn, oHalted);
  not g629 (n_855, \Nanod[permStart] );
  CDN_flop oReset_reg(.clk (clk), .d (n_712), .sena (enT1), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (oReset));
  CDN_flop oHalted_reg(.clk (clk), .d (n_711), .sena (enT1), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (oHalted));
  CDN_flop \rFC_reg[0] (.clk (clk), .d (n_668), .sena (n_667), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q (FC0));
  CDN_flop \rFC_reg[1] (.clk (clk), .d (n_669), .sena (n_667), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q (FC1));
  CDN_flop \rFC_reg[2] (.clk (clk), .d (pswS), .sena (n_667), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q (FC2));
  not g641 (n_868, iplComp);
  CDN_flop intPend_reg(.clk (clk), .d (n_682), .sena (n_876), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (intPend));
  CDN_flop Spuria_reg(.clk (clk), .d (n_877), .sena (enT4), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Spuria));
  CDN_flop Avia_reg(.clk (clk), .d (n_878), .sena (enT4), .aclr (1'b0),
       .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (Avia));
  CDN_flop \inl_reg[0] (.clk (clk), .d (iIpl[0]), .sena (n_880), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b1), .q (inl[0]));
  CDN_flop \inl_reg[1] (.clk (clk), .d (iIpl[1]), .sena (n_880), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b1), .q (inl[1]));
  CDN_flop \inl_reg[2] (.clk (clk), .d (iIpl[2]), .sena (n_880), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b1), .q (inl[2]));
  CDN_flop updIll_reg(.clk (clk), .d (microLatch[0]), .sena (enT4),
       .aclr (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (updIll));
  CDN_flop prevNmi_reg(.clk (clk), .d (nmi), .sena (enPhi2), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (prevNmi));
  CDN_flop E_reg(.clk (clk), .d (n_897), .sena (n_898), .aclr (1'b0),
       .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (E));
  CDN_flop \eCntr_reg[0] (.clk (clk), .d (n_900), .sena (n_901), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (eCntr[0]));
  CDN_flop \eCntr_reg[1] (.clk (clk), .d (n_902), .sena (n_901), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (eCntr[1]));
  CDN_flop \eCntr_reg[2] (.clk (clk), .d (n_903), .sena (n_901), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (eCntr[2]));
  CDN_flop \eCntr_reg[3] (.clk (clk), .d (n_904), .sena (n_901), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (eCntr[3]));
  CDN_flop rVma_reg(.clk (clk), .d (1'b1), .sena (pwrUp), .aclr (1'b0),
       .apre (1'b0), .srl (n_1654), .srd (n_905), .q (VMAn));
  or g661 (n_1654, n_693, n_906);
  CDN_flop iStop_reg(.clk (clk), .d (n_695), .sena (n_918), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q (iStop));
  CDN_flop A0Err_reg(.clk (clk), .d (1'b1), .sena (n_677), .aclr
       (1'b0), .apre (1'b0), .srl (n_1663), .srd (extReset), .q
       (A0Err));
  or g667 (n_1663, n_920, extReset);
  CDN_flop excRst_reg(.clk (clk), .d (1'b0), .sena (1'b0), .aclr
       (1'b0), .apre (1'b0), .srl (n_1669), .srd (extReset), .q
       (excRst));
  or g670 (n_1669, n_921, extReset);
  CDN_flop BerrA_reg(.clk (clk), .d (n_672), .sena (n_925), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q (BerrA));
  CDN_flop rAddrErr_reg(.clk (clk), .d (n_603), .sena (n_929), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (rAddrErr));
  CDN_flop iBusErr_reg(.clk (clk), .d (n_673), .sena (enPhi1), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (iBusErr));
  CDN_flop Err6591_reg(.clk (clk), .d (enErrClk), .sena (enPhi1), .aclr
       (1'b0), .apre (1'b0), .srl (extReset), .srd (1'b0), .q
       (Err6591));
  not g681 (n_930, irdToCcr_t4);
  CDN_flop Tpend_reg(.clk (clk), .d (n_679), .sena (n_935), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (Tpend));
  CDN_flop pswT_reg(.clk (clk), .d (n_716), .sena (n_940), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (pswT));
  CDN_flop pswS_reg(.clk (clk), .d (n_666), .sena (n_940), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (pswS));
  CDN_flop \pswI_reg[0] (.clk (clk), .d (n_713), .sena (n_948), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (pswI[0]));
  CDN_flop \pswI_reg[1] (.clk (clk), .d (n_714), .sena (n_948), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (pswI[1]));
  CDN_flop \pswI_reg[2] (.clk (clk), .d (n_715), .sena (n_948), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (pswI[2]));
  CDN_flop irdToCcr_t4_reg(.clk (clk), .d (\Irdecod[toCcr] ), .sena
       (enT4), .aclr (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0),
       .q (irdToCcr_t4));
  CDN_flop \ftu_reg[0] (.clk (clk), .d (n_650), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[0]));
  CDN_flop \ftu_reg[1] (.clk (clk), .d (n_651), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[1]));
  CDN_flop \ftu_reg[2] (.clk (clk), .d (n_652), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[2]));
  CDN_flop \ftu_reg[3] (.clk (clk), .d (n_653), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[3]));
  CDN_flop \ftu_reg[4] (.clk (clk), .d (n_654), .sena (enT3), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[4]));
  CDN_flop \ftu_reg[5] (.clk (clk), .d (n_655), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[5]));
  CDN_flop \ftu_reg[6] (.clk (clk), .d (n_656), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[6]));
  CDN_flop \ftu_reg[7] (.clk (clk), .d (n_657), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[7]));
  CDN_flop \ftu_reg[8] (.clk (clk), .d (n_658), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[8]));
  CDN_flop \ftu_reg[9] (.clk (clk), .d (n_659), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[9]));
  CDN_flop \ftu_reg[10] (.clk (clk), .d (n_660), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[10]));
  CDN_flop \ftu_reg[11] (.clk (clk), .d (n_661), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[11]));
  CDN_flop \ftu_reg[12] (.clk (clk), .d (n_662), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[12]));
  CDN_flop \ftu_reg[13] (.clk (clk), .d (n_663), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[13]));
  CDN_flop \ftu_reg[14] (.clk (clk), .d (n_664), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[14]));
  CDN_flop \ftu_reg[15] (.clk (clk), .d (n_665), .sena (n_955), .aclr
       (1'b0), .apre (1'b0), .srl (pwrUp), .srd (1'b0), .q (ftu[15]));
  CDN_flop \ssw_reg[0] (.clk (clk), .d (FC0), .sena (n_634), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (ssw[0]));
  CDN_flop \ssw_reg[1] (.clk (clk), .d (FC1), .sena (n_634), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (ssw[1]));
  CDN_flop \ssw_reg[2] (.clk (clk), .d (FC2), .sena (n_634), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (ssw[2]));
  CDN_flop \ssw_reg[3] (.clk (clk), .d (inExcept01), .sena (n_634),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (ssw[3]));
  CDN_flop \ssw_reg[4] (.clk (clk), .d (n_956), .sena (n_634), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (ssw[4]));
  CDN_flop \tvnLatch_reg[0] (.clk (clk), .d (tvn[0]), .sena (n_705),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (tvnLatch[0]));
  CDN_flop \tvnLatch_reg[1] (.clk (clk), .d (tvn[1]), .sena (n_705),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (tvnLatch[1]));
  CDN_flop \tvnLatch_reg[2] (.clk (clk), .d (tvn[2]), .sena (n_705),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (tvnLatch[2]));
  CDN_flop \tvnLatch_reg[3] (.clk (clk), .d (tvn[3]), .sena (n_705),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (tvnLatch[3]));
  CDN_flop inExcept01_reg(.clk (clk), .d (n_957), .sena (n_705), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (inExcept01));
  not g733 (n_860, microLatch[16]);
  nand g734 (n_1774, microLatch[15], n_860);
  not g735 (n_854, n_1774);
  nand g738 (n_1777, microLatch[16], n_857);
  not g739 (n_856, n_1777);
  xnor g740 (n_1778, iIpl[0], rIpl[0]);
  xnor g741 (n_1779, iIpl[1], rIpl[1]);
  xnor g742 (n_1780, iIpl[2], rIpl[2]);
  nand g743 (n_1781, n_1778, n_1779, n_1780);
  not g744 (iplStable, n_1781);
  nand g748 (n_866, iIpl[0], iIpl[1], iIpl[2]);
  not g749 (nmi, n_866);
  nand g758 (n_908, FC0, FC1, FC2);
  not g759 (Iac, n_908);
  nand g764 (n_1798, eCntr[0], n_1072, n_1073, eCntr[3]);
  not g765 (n_684, n_1798);
  nand g779 (n_1810, n_1804, n_1072, n_1073, eCntr[3]);
  not g780 (n_886, n_1810);
  nand g785 (n_1815, n_1811, n_1812, tvnLatch[2], tvnLatch[3]);
  not g786 (n_606, n_1815);
  nand g791 (n_1820, tvnLatch[0], n_1812, tvnLatch[2], tvnLatch[3]);
  not g792 (n_607, n_1820);
  nand g797 (n_1825, tvnLatch[0], tvnLatch[1], tvnLatch[2],
       tvnLatch[3]);
  not g798 (n_609, n_1825);
  nor g800 (n_1826, tvn[3], tvn[2], tvn[1]);
  nand g801 (n_957, n_1826, tvn[0]);
  not g802 (n_1804, eCntr[0]);
  not g803 (n_1811, tvnLatch[0]);
  not g804 (n_1812, tvnLatch[1]);
  or g805 (wClk, waitBusCycle, n_881, iAddrErr, Err6591);
  or g806 (n_1829, n_815, n_813);
  or g807 (n_817, n_811, n_809, n_810, n_1829);
  or g808 (n_1830, n_649, \Nanod[abl2Pren] );
  or g809 (n_1831, \Nanod[const2Ftu] , \Nanod[pswIToFtu] );
  or g810 (n_1832, \Nanod[ird2Ftu] , \Nanod[sr2Ftu] );
  or g811 (n_954, \Nanod[tvn2Ftu] , n_1830, n_1831, n_1832);
  nor g812 (n_1833, eCntr[3], eCntr[2]);
  and g813 (n_1834, enPhi2, addrOe);
  and g814 (n_1835, n_872, eCntr[0]);
  and g815 (n_693, eCntr[1], n_1833, n_1834, n_1835);
  nor g816 (n_1837, eCntr[3], eCntr[2]);
  and g817 (n_1838, n_1836, enPhi1);
  not g818 (n_1836, eCntr[1]);
  and g819 (n_906, n_1804, n_905, n_1837, n_1838);
  and g820 (n_869, inl[0], inl[1], inl[2], Iac);
endmodule

`ifdef RC_CDN_GENERIC_GATE
`else
module CDN_dc(cf, dcf, z);
  input cf, dcf;
  output z;
  wire cf, dcf;
  wire z;
  assign z = dcf ? 1'bx : cf;
endmodule
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
module CDN_flop(clk, d, sena, aclr, apre, srl, srd, q);
  input clk, d, sena, aclr, apre, srl, srd;
  output q;
  wire clk, d, sena, aclr, apre, srl, srd;
  wire q;
  reg  qi;
  assign #1 q = qi;
  always 
    @(posedge clk or posedge apre or posedge aclr) 
      if (aclr) 
        qi <= 0;
      else if (apre) 
          qi <= 1;
        else if (srl) 
            qi <= srd;
          else begin
            if (sena) 
              qi <= d;
          end
  initial 
    qi <= 1'b0;
endmodule
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux136(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, sel13,
     data13, sel14, data14, sel15, data15, sel16, data16, sel17,
     data17, sel18, data18, sel19, data19, sel20, data20, sel21,
     data21, sel22, data22, sel23, data23, sel24, data24, sel25,
     data25, sel26, data26, sel27, data27, sel28, data28, sel29,
     data29, sel30, data30, sel31, data31, sel32, data32, sel33,
     data33, sel34, data34, sel35, data35, sel36, data36, sel37,
     data37, sel38, data38, sel39, data39, sel40, data40, sel41,
     data41, sel42, data42, sel43, data43, sel44, data44, sel45,
     data45, sel46, data46, sel47, data47, sel48, data48, sel49,
     data49, sel50, data50, sel51, data51, sel52, data52, sel53,
     data53, sel54, data54, sel55, data55, sel56, data56, sel57,
     data57, sel58, data58, sel59, data59, sel60, data60, sel61,
     data61, sel62, data62, sel63, data63, sel64, data64, sel65,
     data65, sel66, data66, sel67, data67, sel68, data68, sel69,
     data69, sel70, data70, sel71, data71, sel72, data72, sel73,
     data73, sel74, data74, sel75, data75, sel76, data76, sel77,
     data77, sel78, data78, sel79, data79, sel80, data80, sel81,
     data81, sel82, data82, sel83, data83, sel84, data84, sel85,
     data85, sel86, data86, sel87, data87, sel88, data88, sel89,
     data89, sel90, data90, sel91, data91, sel92, data92, sel93,
     data93, sel94, data94, sel95, data95, sel96, data96, sel97,
     data97, sel98, data98, sel99, data99, sel100, data100, sel101,
     data101, sel102, data102, sel103, data103, sel104, data104,
     sel105, data105, sel106, data106, sel107, data107, sel108,
     data108, sel109, data109, sel110, data110, sel111, data111,
     sel112, data112, sel113, data113, sel114, data114, sel115,
     data115, sel116, data116, sel117, data117, sel118, data118,
     sel119, data119, sel120, data120, sel121, data121, sel122,
     data122, sel123, data123, sel124, data124, sel125, data125,
     sel126, data126, sel127, data127, sel128, data128, sel129,
     data129, sel130, data130, sel131, data131, sel132, data132,
     sel133, data133, sel134, data134, sel135, data135, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12, sel13,
       data13, sel14, data14, sel15, data15, sel16, data16, sel17,
       data17, sel18, data18, sel19, data19, sel20, data20, sel21,
       data21, sel22, data22, sel23, data23, sel24, data24, sel25,
       data25, sel26, data26, sel27, data27, sel28, data28, sel29,
       data29, sel30, data30, sel31, data31, sel32, data32, sel33,
       data33, sel34, data34, sel35, data35, sel36, data36, sel37,
       data37, sel38, data38, sel39, data39, sel40, data40, sel41,
       data41, sel42, data42, sel43, data43, sel44, data44, sel45,
       data45, sel46, data46, sel47, data47, sel48, data48, sel49,
       data49, sel50, data50, sel51, data51, sel52, data52, sel53,
       data53, sel54, data54, sel55, data55, sel56, data56, sel57,
       data57, sel58, data58, sel59, data59, sel60, data60, sel61,
       data61, sel62, data62, sel63, data63, sel64, data64, sel65,
       data65, sel66, data66, sel67, data67, sel68, data68, sel69,
       data69, sel70, data70, sel71, data71, sel72, data72, sel73,
       data73, sel74, data74, sel75, data75, sel76, data76, sel77,
       data77, sel78, data78, sel79, data79, sel80, data80, sel81,
       data81, sel82, data82, sel83, data83, sel84, data84, sel85,
       data85, sel86, data86, sel87, data87, sel88, data88, sel89,
       data89, sel90, data90, sel91, data91, sel92, data92, sel93,
       data93, sel94, data94, sel95, data95, sel96, data96, sel97,
       data97, sel98, data98, sel99, data99, sel100, data100, sel101,
       data101, sel102, data102, sel103, data103, sel104, data104,
       sel105, data105, sel106, data106, sel107, data107, sel108,
       data108, sel109, data109, sel110, data110, sel111, data111,
       sel112, data112, sel113, data113, sel114, data114, sel115,
       data115, sel116, data116, sel117, data117, sel118, data118,
       sel119, data119, sel120, data120, sel121, data121, sel122,
       data122, sel123, data123, sel124, data124, sel125, data125,
       sel126, data126, sel127, data127, sel128, data128, sel129,
       data129, sel130, data130, sel131, data131, sel132, data132,
       sel133, data133, sel134, data134, sel135, data135;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12, sel13, data13,
       sel14, data14, sel15, data15, sel16, data16, sel17, data17,
       sel18, data18, sel19, data19, sel20, data20, sel21, data21,
       sel22, data22, sel23, data23, sel24, data24, sel25, data25,
       sel26, data26, sel27, data27, sel28, data28, sel29, data29,
       sel30, data30, sel31, data31, sel32, data32, sel33, data33,
       sel34, data34, sel35, data35, sel36, data36, sel37, data37,
       sel38, data38, sel39, data39, sel40, data40, sel41, data41,
       sel42, data42, sel43, data43, sel44, data44, sel45, data45,
       sel46, data46, sel47, data47, sel48, data48, sel49, data49,
       sel50, data50, sel51, data51, sel52, data52, sel53, data53,
       sel54, data54, sel55, data55, sel56, data56, sel57, data57,
       sel58, data58, sel59, data59, sel60, data60, sel61, data61,
       sel62, data62, sel63, data63, sel64, data64, sel65, data65,
       sel66, data66, sel67, data67, sel68, data68, sel69, data69,
       sel70, data70, sel71, data71, sel72, data72, sel73, data73,
       sel74, data74, sel75, data75, sel76, data76, sel77, data77,
       sel78, data78, sel79, data79, sel80, data80, sel81, data81,
       sel82, data82, sel83, data83, sel84, data84, sel85, data85,
       sel86, data86, sel87, data87, sel88, data88, sel89, data89,
       sel90, data90, sel91, data91, sel92, data92, sel93, data93,
       sel94, data94, sel95, data95, sel96, data96, sel97, data97,
       sel98, data98, sel99, data99, sel100, data100, sel101, data101,
       sel102, data102, sel103, data103, sel104, data104, sel105,
       data105, sel106, data106, sel107, data107, sel108, data108,
       sel109, data109, sel110, data110, sel111, data111, sel112,
       data112, sel113, data113, sel114, data114, sel115, data115,
       sel116, data116, sel117, data117, sel118, data118, sel119,
       data119, sel120, data120, sel121, data121, sel122, data122,
       sel123, data123, sel124, data124, sel125, data125, sel126,
       data126, sel127, data127, sel128, data128, sel129, data129,
       sel130, data130, sel131, data131, sel132, data132, sel133,
       data133, sel134, data134, sel135, data135;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or sel9 or sel10 or sel11 or sel12 or sel13 or sel14 or
         sel15 or sel16 or sel17 or sel18 or sel19 or sel20 or sel21 or
         sel22 or sel23 or sel24 or sel25 or sel26 or sel27 or sel28 or
         sel29 or sel30 or sel31 or sel32 or sel33 or sel34 or sel35 or
         sel36 or sel37 or sel38 or sel39 or sel40 or sel41 or sel42 or
         sel43 or sel44 or sel45 or sel46 or sel47 or sel48 or sel49 or
         sel50 or sel51 or sel52 or sel53 or sel54 or sel55 or sel56 or
         sel57 or sel58 or sel59 or sel60 or sel61 or sel62 or sel63 or
         sel64 or sel65 or sel66 or sel67 or sel68 or sel69 or sel70 or
         sel71 or sel72 or sel73 or sel74 or sel75 or sel76 or sel77 or
         sel78 or sel79 or sel80 or sel81 or sel82 or sel83 or sel84 or
         sel85 or sel86 or sel87 or sel88 or sel89 or sel90 or sel91 or
         sel92 or sel93 or sel94 or sel95 or sel96 or sel97 or sel98 or
         sel99 or sel100 or sel101 or sel102 or sel103 or sel104 or
         sel105 or sel106 or sel107 or sel108 or sel109 or sel110 or
         sel111 or sel112 or sel113 or sel114 or sel115 or sel116 or
         sel117 or sel118 or sel119 or sel120 or sel121 or sel122 or
         sel123 or sel124 or sel125 or sel126 or sel127 or sel128 or
         sel129 or sel130 or sel131 or sel132 or sel133 or sel134 or
         sel135 or data0 or data1 or data2 or data3 or data4 or data5
         or data6 or data7 or data8 or data9 or data10 or data11 or
         data12 or data13 or data14 or data15 or data16 or data17 or
         data18 or data19 or data20 or data21 or data22 or data23 or
         data24 or data25 or data26 or data27 or data28 or data29 or
         data30 or data31 or data32 or data33 or data34 or data35 or
         data36 or data37 or data38 or data39 or data40 or data41 or
         data42 or data43 or data44 or data45 or data46 or data47 or
         data48 or data49 or data50 or data51 or data52 or data53 or
         data54 or data55 or data56 or data57 or data58 or data59 or
         data60 or data61 or data62 or data63 or data64 or data65 or
         data66 or data67 or data68 or data69 or data70 or data71 or
         data72 or data73 or data74 or data75 or data76 or data77 or
         data78 or data79 or data80 or data81 or data82 or data83 or
         data84 or data85 or data86 or data87 or data88 or data89 or
         data90 or data91 or data92 or data93 or data94 or data95 or
         data96 or data97 or data98 or data99 or data100 or data101 or
         data102 or data103 or data104 or data105 or data106 or data107
         or data108 or data109 or data110 or data111 or data112 or
         data113 or data114 or data115 or data116 or data117 or data118
         or data119 or data120 or data121 or data122 or data123 or
         data124 or data125 or data126 or data127 or data128 or data129
         or data130 or data131 or data132 or data133 or data134 or
         data135) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
           sel9, sel10, sel11, sel12, sel13, sel14, sel15, sel16,
           sel17, sel18, sel19, sel20, sel21, sel22, sel23, sel24,
           sel25, sel26, sel27, sel28, sel29, sel30, sel31, sel32,
           sel33, sel34, sel35, sel36, sel37, sel38, sel39, sel40,
           sel41, sel42, sel43, sel44, sel45, sel46, sel47, sel48,
           sel49, sel50, sel51, sel52, sel53, sel54, sel55, sel56,
           sel57, sel58, sel59, sel60, sel61, sel62, sel63, sel64,
           sel65, sel66, sel67, sel68, sel69, sel70, sel71, sel72,
           sel73, sel74, sel75, sel76, sel77, sel78, sel79, sel80,
           sel81, sel82, sel83, sel84, sel85, sel86, sel87, sel88,
           sel89, sel90, sel91, sel92, sel93, sel94, sel95, sel96,
           sel97, sel98, sel99, sel100, sel101, sel102, sel103, sel104,
           sel105, sel106, sel107, sel108, sel109, sel110, sel111,
           sel112, sel113, sel114, sel115, sel116, sel117, sel118,
           sel119, sel120, sel121, sel122, sel123, sel124, sel125,
           sel126, sel127, sel128, sel129, sel130, sel131, sel132,
           sel133, sel134, sel135})
       136'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data0;
       136'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data1;
       136'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data2;
       136'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data3;
       136'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data4;
       136'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data5;
       136'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data6;
       136'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data7;
       136'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data8;
       136'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data9;
       136'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data10;
       136'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data11;
       136'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data12;
       136'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data13;
       136'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data14;
       136'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data15;
       136'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data16;
       136'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data17;
       136'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data18;
       136'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data19;
       136'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data20;
       136'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data21;
       136'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data22;
       136'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data23;
       136'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data24;
       136'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data25;
       136'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data26;
       136'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data27;
       136'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data28;
       136'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data29;
       136'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data30;
       136'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data31;
       136'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data32;
       136'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data33;
       136'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data34;
       136'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data35;
       136'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data36;
       136'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data37;
       136'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data38;
       136'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data39;
       136'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data40;
       136'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data41;
       136'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data42;
       136'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data43;
       136'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data44;
       136'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data45;
       136'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data46;
       136'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data47;
       136'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data48;
       136'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data49;
       136'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data50;
       136'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data51;
       136'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data52;
       136'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data53;
       136'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data54;
       136'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data55;
       136'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data56;
       136'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data57;
       136'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data58;
       136'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data59;
       136'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data60;
       136'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data61;
       136'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data62;
       136'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000:
           z = data63;
       136'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000:
           z = data64;
       136'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000:
           z = data65;
       136'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000:
           z = data66;
       136'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000:
           z = data67;
       136'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000:
           z = data68;
       136'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000:
           z = data69;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000:
           z = data70;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000:
           z = data71;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000:
           z = data72;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000:
           z = data73;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000:
           z = data74;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000:
           z = data75;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000:
           z = data76;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000:
           z = data77;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000:
           z = data78;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000:
           z = data79;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000:
           z = data80;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000:
           z = data81;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000:
           z = data82;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000:
           z = data83;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000:
           z = data84;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000:
           z = data85;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000:
           z = data86;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000:
           z = data87;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000:
           z = data88;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000:
           z = data89;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000:
           z = data90;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000:
           z = data91;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000:
           z = data92;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000:
           z = data93;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000:
           z = data94;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000:
           z = data95;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000:
           z = data96;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000:
           z = data97;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000:
           z = data98;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000:
           z = data99;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000:
           z = data100;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000:
           z = data101;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000:
           z = data102;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000:
           z = data103;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000:
           z = data104;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000:
           z = data105;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000:
           z = data106;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000:
           z = data107;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000:
           z = data108;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000:
           z = data109;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000:
           z = data110;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000:
           z = data111;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000:
           z = data112;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000:
           z = data113;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000:
           z = data114;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000:
           z = data115;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000:
           z = data116;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000:
           z = data117;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000:
           z = data118;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000:
           z = data119;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000:
           z = data120;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000:
           z = data121;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000:
           z = data122;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000:
           z = data123;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000:
           z = data124;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000:
           z = data125;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000:
           z = data126;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000:
           z = data127;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000:
           z = data128;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000:
           z = data129;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000:
           z = data130;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000:
           z = data131;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000:
           z = data132;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100:
           z = data133;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010:
           z = data134;
       136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001:
           z = data135;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux136(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, sel13,
     data13, sel14, data14, sel15, data15, sel16, data16, sel17,
     data17, sel18, data18, sel19, data19, sel20, data20, sel21,
     data21, sel22, data22, sel23, data23, sel24, data24, sel25,
     data25, sel26, data26, sel27, data27, sel28, data28, sel29,
     data29, sel30, data30, sel31, data31, sel32, data32, sel33,
     data33, sel34, data34, sel35, data35, sel36, data36, sel37,
     data37, sel38, data38, sel39, data39, sel40, data40, sel41,
     data41, sel42, data42, sel43, data43, sel44, data44, sel45,
     data45, sel46, data46, sel47, data47, sel48, data48, sel49,
     data49, sel50, data50, sel51, data51, sel52, data52, sel53,
     data53, sel54, data54, sel55, data55, sel56, data56, sel57,
     data57, sel58, data58, sel59, data59, sel60, data60, sel61,
     data61, sel62, data62, sel63, data63, sel64, data64, sel65,
     data65, sel66, data66, sel67, data67, sel68, data68, sel69,
     data69, sel70, data70, sel71, data71, sel72, data72, sel73,
     data73, sel74, data74, sel75, data75, sel76, data76, sel77,
     data77, sel78, data78, sel79, data79, sel80, data80, sel81,
     data81, sel82, data82, sel83, data83, sel84, data84, sel85,
     data85, sel86, data86, sel87, data87, sel88, data88, sel89,
     data89, sel90, data90, sel91, data91, sel92, data92, sel93,
     data93, sel94, data94, sel95, data95, sel96, data96, sel97,
     data97, sel98, data98, sel99, data99, sel100, data100, sel101,
     data101, sel102, data102, sel103, data103, sel104, data104,
     sel105, data105, sel106, data106, sel107, data107, sel108,
     data108, sel109, data109, sel110, data110, sel111, data111,
     sel112, data112, sel113, data113, sel114, data114, sel115,
     data115, sel116, data116, sel117, data117, sel118, data118,
     sel119, data119, sel120, data120, sel121, data121, sel122,
     data122, sel123, data123, sel124, data124, sel125, data125,
     sel126, data126, sel127, data127, sel128, data128, sel129,
     data129, sel130, data130, sel131, data131, sel132, data132,
     sel133, data133, sel134, data134, sel135, data135, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12, sel13,
       data13, sel14, data14, sel15, data15, sel16, data16, sel17,
       data17, sel18, data18, sel19, data19, sel20, data20, sel21,
       data21, sel22, data22, sel23, data23, sel24, data24, sel25,
       data25, sel26, data26, sel27, data27, sel28, data28, sel29,
       data29, sel30, data30, sel31, data31, sel32, data32, sel33,
       data33, sel34, data34, sel35, data35, sel36, data36, sel37,
       data37, sel38, data38, sel39, data39, sel40, data40, sel41,
       data41, sel42, data42, sel43, data43, sel44, data44, sel45,
       data45, sel46, data46, sel47, data47, sel48, data48, sel49,
       data49, sel50, data50, sel51, data51, sel52, data52, sel53,
       data53, sel54, data54, sel55, data55, sel56, data56, sel57,
       data57, sel58, data58, sel59, data59, sel60, data60, sel61,
       data61, sel62, data62, sel63, data63, sel64, data64, sel65,
       data65, sel66, data66, sel67, data67, sel68, data68, sel69,
       data69, sel70, data70, sel71, data71, sel72, data72, sel73,
       data73, sel74, data74, sel75, data75, sel76, data76, sel77,
       data77, sel78, data78, sel79, data79, sel80, data80, sel81,
       data81, sel82, data82, sel83, data83, sel84, data84, sel85,
       data85, sel86, data86, sel87, data87, sel88, data88, sel89,
       data89, sel90, data90, sel91, data91, sel92, data92, sel93,
       data93, sel94, data94, sel95, data95, sel96, data96, sel97,
       data97, sel98, data98, sel99, data99, sel100, data100, sel101,
       data101, sel102, data102, sel103, data103, sel104, data104,
       sel105, data105, sel106, data106, sel107, data107, sel108,
       data108, sel109, data109, sel110, data110, sel111, data111,
       sel112, data112, sel113, data113, sel114, data114, sel115,
       data115, sel116, data116, sel117, data117, sel118, data118,
       sel119, data119, sel120, data120, sel121, data121, sel122,
       data122, sel123, data123, sel124, data124, sel125, data125,
       sel126, data126, sel127, data127, sel128, data128, sel129,
       data129, sel130, data130, sel131, data131, sel132, data132,
       sel133, data133, sel134, data134, sel135, data135;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12, sel13, data13,
       sel14, data14, sel15, data15, sel16, data16, sel17, data17,
       sel18, data18, sel19, data19, sel20, data20, sel21, data21,
       sel22, data22, sel23, data23, sel24, data24, sel25, data25,
       sel26, data26, sel27, data27, sel28, data28, sel29, data29,
       sel30, data30, sel31, data31, sel32, data32, sel33, data33,
       sel34, data34, sel35, data35, sel36, data36, sel37, data37,
       sel38, data38, sel39, data39, sel40, data40, sel41, data41,
       sel42, data42, sel43, data43, sel44, data44, sel45, data45,
       sel46, data46, sel47, data47, sel48, data48, sel49, data49,
       sel50, data50, sel51, data51, sel52, data52, sel53, data53,
       sel54, data54, sel55, data55, sel56, data56, sel57, data57,
       sel58, data58, sel59, data59, sel60, data60, sel61, data61,
       sel62, data62, sel63, data63, sel64, data64, sel65, data65,
       sel66, data66, sel67, data67, sel68, data68, sel69, data69,
       sel70, data70, sel71, data71, sel72, data72, sel73, data73,
       sel74, data74, sel75, data75, sel76, data76, sel77, data77,
       sel78, data78, sel79, data79, sel80, data80, sel81, data81,
       sel82, data82, sel83, data83, sel84, data84, sel85, data85,
       sel86, data86, sel87, data87, sel88, data88, sel89, data89,
       sel90, data90, sel91, data91, sel92, data92, sel93, data93,
       sel94, data94, sel95, data95, sel96, data96, sel97, data97,
       sel98, data98, sel99, data99, sel100, data100, sel101, data101,
       sel102, data102, sel103, data103, sel104, data104, sel105,
       data105, sel106, data106, sel107, data107, sel108, data108,
       sel109, data109, sel110, data110, sel111, data111, sel112,
       data112, sel113, data113, sel114, data114, sel115, data115,
       sel116, data116, sel117, data117, sel118, data118, sel119,
       data119, sel120, data120, sel121, data121, sel122, data122,
       sel123, data123, sel124, data124, sel125, data125, sel126,
       data126, sel127, data127, sel128, data128, sel129, data129,
       sel130, data130, sel131, data131, sel132, data132, sel133,
       data133, sel134, data134, sel135, data135;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8, w_9, w_10, w_11, w_12, w_13, w_14, w_15;
  wire w_16, w_17, w_18, w_19, w_20, w_21, w_22, w_23;
  wire w_24, w_25, w_26, w_27, w_28, w_29, w_30, w_31;
  wire w_32, w_33, w_34, w_35, w_36, w_37, w_38, w_39;
  wire w_40, w_41, w_42, w_43, w_44, w_45, w_46, w_47;
  wire w_48, w_49, w_50, w_51, w_52, w_53, w_54, w_55;
  wire w_56, w_57, w_58, w_59, w_60, w_61, w_62, w_63;
  wire w_64, w_65, w_66, w_67, w_68, w_69, w_70, w_71;
  wire w_72, w_73, w_74, w_75, w_76, w_77, w_78, w_79;
  wire w_80, w_81, w_82, w_83, w_84, w_85, w_86, w_87;
  wire w_88, w_89, w_90, w_91, w_92, w_93, w_94, w_95;
  wire w_96, w_97, w_98, w_99, w_100, w_101, w_102, w_103;
  wire w_104, w_105, w_106, w_107, w_108, w_109, w_110, w_111;
  wire w_112, w_113, w_114, w_115, w_116, w_117, w_118, w_119;
  wire w_120, w_121, w_122, w_123, w_124, w_125, w_126, w_127;
  wire w_128, w_129, w_130, w_131, w_132, w_133, w_134, w_135;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  and a_9 (w_9, sel9, data9);
  and a_10 (w_10, sel10, data10);
  and a_11 (w_11, sel11, data11);
  and a_12 (w_12, sel12, data12);
  and a_13 (w_13, sel13, data13);
  and a_14 (w_14, sel14, data14);
  and a_15 (w_15, sel15, data15);
  and a_16 (w_16, sel16, data16);
  and a_17 (w_17, sel17, data17);
  and a_18 (w_18, sel18, data18);
  and a_19 (w_19, sel19, data19);
  and a_20 (w_20, sel20, data20);
  and a_21 (w_21, sel21, data21);
  and a_22 (w_22, sel22, data22);
  and a_23 (w_23, sel23, data23);
  and a_24 (w_24, sel24, data24);
  and a_25 (w_25, sel25, data25);
  and a_26 (w_26, sel26, data26);
  and a_27 (w_27, sel27, data27);
  and a_28 (w_28, sel28, data28);
  and a_29 (w_29, sel29, data29);
  and a_30 (w_30, sel30, data30);
  and a_31 (w_31, sel31, data31);
  and a_32 (w_32, sel32, data32);
  and a_33 (w_33, sel33, data33);
  and a_34 (w_34, sel34, data34);
  and a_35 (w_35, sel35, data35);
  and a_36 (w_36, sel36, data36);
  and a_37 (w_37, sel37, data37);
  and a_38 (w_38, sel38, data38);
  and a_39 (w_39, sel39, data39);
  and a_40 (w_40, sel40, data40);
  and a_41 (w_41, sel41, data41);
  and a_42 (w_42, sel42, data42);
  and a_43 (w_43, sel43, data43);
  and a_44 (w_44, sel44, data44);
  and a_45 (w_45, sel45, data45);
  and a_46 (w_46, sel46, data46);
  and a_47 (w_47, sel47, data47);
  and a_48 (w_48, sel48, data48);
  and a_49 (w_49, sel49, data49);
  and a_50 (w_50, sel50, data50);
  and a_51 (w_51, sel51, data51);
  and a_52 (w_52, sel52, data52);
  and a_53 (w_53, sel53, data53);
  and a_54 (w_54, sel54, data54);
  and a_55 (w_55, sel55, data55);
  and a_56 (w_56, sel56, data56);
  and a_57 (w_57, sel57, data57);
  and a_58 (w_58, sel58, data58);
  and a_59 (w_59, sel59, data59);
  and a_60 (w_60, sel60, data60);
  and a_61 (w_61, sel61, data61);
  and a_62 (w_62, sel62, data62);
  and a_63 (w_63, sel63, data63);
  and a_64 (w_64, sel64, data64);
  and a_65 (w_65, sel65, data65);
  and a_66 (w_66, sel66, data66);
  and a_67 (w_67, sel67, data67);
  and a_68 (w_68, sel68, data68);
  and a_69 (w_69, sel69, data69);
  and a_70 (w_70, sel70, data70);
  and a_71 (w_71, sel71, data71);
  and a_72 (w_72, sel72, data72);
  and a_73 (w_73, sel73, data73);
  and a_74 (w_74, sel74, data74);
  and a_75 (w_75, sel75, data75);
  and a_76 (w_76, sel76, data76);
  and a_77 (w_77, sel77, data77);
  and a_78 (w_78, sel78, data78);
  and a_79 (w_79, sel79, data79);
  and a_80 (w_80, sel80, data80);
  and a_81 (w_81, sel81, data81);
  and a_82 (w_82, sel82, data82);
  and a_83 (w_83, sel83, data83);
  and a_84 (w_84, sel84, data84);
  and a_85 (w_85, sel85, data85);
  and a_86 (w_86, sel86, data86);
  and a_87 (w_87, sel87, data87);
  and a_88 (w_88, sel88, data88);
  and a_89 (w_89, sel89, data89);
  and a_90 (w_90, sel90, data90);
  and a_91 (w_91, sel91, data91);
  and a_92 (w_92, sel92, data92);
  and a_93 (w_93, sel93, data93);
  and a_94 (w_94, sel94, data94);
  and a_95 (w_95, sel95, data95);
  and a_96 (w_96, sel96, data96);
  and a_97 (w_97, sel97, data97);
  and a_98 (w_98, sel98, data98);
  and a_99 (w_99, sel99, data99);
  and a_100 (w_100, sel100, data100);
  and a_101 (w_101, sel101, data101);
  and a_102 (w_102, sel102, data102);
  and a_103 (w_103, sel103, data103);
  and a_104 (w_104, sel104, data104);
  and a_105 (w_105, sel105, data105);
  and a_106 (w_106, sel106, data106);
  and a_107 (w_107, sel107, data107);
  and a_108 (w_108, sel108, data108);
  and a_109 (w_109, sel109, data109);
  and a_110 (w_110, sel110, data110);
  and a_111 (w_111, sel111, data111);
  and a_112 (w_112, sel112, data112);
  and a_113 (w_113, sel113, data113);
  and a_114 (w_114, sel114, data114);
  and a_115 (w_115, sel115, data115);
  and a_116 (w_116, sel116, data116);
  and a_117 (w_117, sel117, data117);
  and a_118 (w_118, sel118, data118);
  and a_119 (w_119, sel119, data119);
  and a_120 (w_120, sel120, data120);
  and a_121 (w_121, sel121, data121);
  and a_122 (w_122, sel122, data122);
  and a_123 (w_123, sel123, data123);
  and a_124 (w_124, sel124, data124);
  and a_125 (w_125, sel125, data125);
  and a_126 (w_126, sel126, data126);
  and a_127 (w_127, sel127, data127);
  and a_128 (w_128, sel128, data128);
  and a_129 (w_129, sel129, data129);
  and a_130 (w_130, sel130, data130);
  and a_131 (w_131, sel131, data131);
  and a_132 (w_132, sel132, data132);
  and a_133 (w_133, sel133, data133);
  and a_134 (w_134, sel134, data134);
  and a_135 (w_135, sel135, data135);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11, w_12, w_13, w_14, w_15, w_16, w_17, w_18, w_19, w_20,
       w_21, w_22, w_23, w_24, w_25, w_26, w_27, w_28, w_29, w_30,
       w_31, w_32, w_33, w_34, w_35, w_36, w_37, w_38, w_39, w_40,
       w_41, w_42, w_43, w_44, w_45, w_46, w_47, w_48, w_49, w_50,
       w_51, w_52, w_53, w_54, w_55, w_56, w_57, w_58, w_59, w_60,
       w_61, w_62, w_63, w_64, w_65, w_66, w_67, w_68, w_69, w_70,
       w_71, w_72, w_73, w_74, w_75, w_76, w_77, w_78, w_79, w_80,
       w_81, w_82, w_83, w_84, w_85, w_86, w_87, w_88, w_89, w_90,
       w_91, w_92, w_93, w_94, w_95, w_96, w_97, w_98, w_99, w_100,
       w_101, w_102, w_103, w_104, w_105, w_106, w_107, w_108, w_109,
       w_110, w_111, w_112, w_113, w_114, w_115, w_116, w_117, w_118,
       w_119, w_120, w_121, w_122, w_123, w_124, w_125, w_126, w_127,
       w_128, w_129, w_130, w_131, w_132, w_133, w_134, w_135);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux9(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or data0 or data1 or data2 or data3 or data4 or data5 or
         data6 or data7 or data8) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8})
       9'b100000000: z = data0;
       9'b010000000: z = data1;
       9'b001000000: z = data2;
       9'b000100000: z = data3;
       9'b000010000: z = data4;
       9'b000001000: z = data5;
       9'b000000100: z = data6;
       9'b000000010: z = data7;
       9'b000000001: z = data8;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux9(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux8(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         data0 or data1 or data2 or data3 or data4 or data5 or data6 or
         data7) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7})
       8'b10000000: z = data0;
       8'b01000000: z = data1;
       8'b00100000: z = data2;
       8'b00010000: z = data3;
       8'b00001000: z = data4;
       8'b00000100: z = data5;
       8'b00000010: z = data6;
       8'b00000001: z = data7;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux8(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux12(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or sel9 or sel10 or sel11 or data0 or data1 or data2 or
         data3 or data4 or data5 or data6 or data7 or data8 or data9 or
         data10 or data11) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
           sel9, sel10, sel11})
       12'b100000000000: z = data0;
       12'b010000000000: z = data1;
       12'b001000000000: z = data2;
       12'b000100000000: z = data3;
       12'b000010000000: z = data4;
       12'b000001000000: z = data5;
       12'b000000100000: z = data6;
       12'b000000010000: z = data7;
       12'b000000001000: z = data8;
       12'b000000000100: z = data9;
       12'b000000000010: z = data10;
       12'b000000000001: z = data11;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux12(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8, w_9, w_10, w_11;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  and a_9 (w_9, sel9, data9);
  and a_10 (w_10, sel10, data10);
  and a_11 (w_11, sel11, data11);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux10(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or sel9 or data0 or data1 or data2 or data3 or data4 or
         data5 or data6 or data7 or data8 or data9) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
           sel9})
       10'b1000000000: z = data0;
       10'b0100000000: z = data1;
       10'b0010000000: z = data2;
       10'b0001000000: z = data3;
       10'b0000100000: z = data4;
       10'b0000010000: z = data5;
       10'b0000001000: z = data6;
       10'b0000000100: z = data7;
       10'b0000000010: z = data8;
       10'b0000000001: z = data9;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux10(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8, w_9;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  and a_9 (w_9, sel9, data9);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux7(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or data0 or
         data1 or data2 or data3 or data4 or data5 or data6) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6})
       7'b1000000: z = data0;
       7'b0100000: z = data1;
       7'b0010000: z = data2;
       7'b0001000: z = data3;
       7'b0000100: z = data4;
       7'b0000010: z = data5;
       7'b0000001: z = data6;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux7(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux5(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or data0 or data1 or data2
         or data3 or data4) 
      case ({sel0, sel1, sel2, sel3, sel4})
       5'b10000: z = data0;
       5'b01000: z = data1;
       5'b00100: z = data2;
       5'b00010: z = data3;
       5'b00001: z = data4;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux5(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  or org (z, w_0, w_1, w_2, w_3, w_4);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux2(sel0, data0, sel1, data1, z);
  input sel0, data0, sel1, data1;
  output z;
  wire sel0, data0, sel1, data1;
  reg  z;
  always 
    @(sel0 or sel1 or data0 or data1) 
      case ({sel0, sel1})
       2'b10: z = data0;
       2'b01: z = data1;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux2(sel0, data0, sel1, data1, z);
  input sel0, data0, sel1, data1;
  output z;
  wire sel0, data0, sel1, data1;
  wire z;
  wire w_0, w_1;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  or org (z, w_0, w_1);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux11(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or sel9 or sel10 or data0 or data1 or data2 or data3 or
         data4 or data5 or data6 or data7 or data8 or data9 or data10) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
           sel9, sel10})
       11'b10000000000: z = data0;
       11'b01000000000: z = data1;
       11'b00100000000: z = data2;
       11'b00010000000: z = data3;
       11'b00001000000: z = data4;
       11'b00000100000: z = data5;
       11'b00000010000: z = data6;
       11'b00000001000: z = data7;
       11'b00000000100: z = data8;
       11'b00000000010: z = data9;
       11'b00000000001: z = data10;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux11(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8, w_9, w_10;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  and a_9 (w_9, sel9, data9);
  and a_10 (w_10, sel10, data10);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux4(sel0, data0, sel1, data1, sel2, data2, sel3, data3, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or data0 or data1 or data2 or data3) 
      case ({sel0, sel1, sel2, sel3})
       4'b1000: z = data0;
       4'b0100: z = data1;
       4'b0010: z = data2;
       4'b0001: z = data3;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux4(sel0, data0, sel1, data1, sel2, data2, sel3, data3, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3;
  wire z;
  wire w_0, w_1, w_2, w_3;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  or org (z, w_0, w_1, w_2, w_3);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux6(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or data0 or data1 or
         data2 or data3 or data4 or data5) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5})
       6'b100000: z = data0;
       6'b010000: z = data1;
       6'b001000: z = data2;
       6'b000100: z = data3;
       6'b000010: z = data4;
       6'b000001: z = data5;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux6(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux3(sel0, data0, sel1, data1, sel2, data2, z);
  input sel0, data0, sel1, data1, sel2, data2;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or data0 or data1 or data2) 
      case ({sel0, sel1, sel2})
       3'b100: z = data0;
       3'b010: z = data1;
       3'b001: z = data2;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux3(sel0, data0, sel1, data1, sel2, data2, z);
  input sel0, data0, sel1, data1, sel2, data2;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2;
  wire z;
  wire w_0, w_1, w_2;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  or org (z, w_0, w_1, w_2);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux13(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or sel9 or sel10 or sel11 or sel12 or data0 or data1 or
         data2 or data3 or data4 or data5 or data6 or data7 or data8 or
         data9 or data10 or data11 or data12) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
           sel9, sel10, sel11, sel12})
       13'b1000000000000: z = data0;
       13'b0100000000000: z = data1;
       13'b0010000000000: z = data2;
       13'b0001000000000: z = data3;
       13'b0000100000000: z = data4;
       13'b0000010000000: z = data5;
       13'b0000001000000: z = data6;
       13'b0000000100000: z = data7;
       13'b0000000010000: z = data8;
       13'b0000000001000: z = data9;
       13'b0000000000100: z = data10;
       13'b0000000000010: z = data11;
       13'b0000000000001: z = data12;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux13(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8, w_9, w_10, w_11, w_12;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  and a_9 (w_9, sel9, data9);
  and a_10 (w_10, sel10, data10);
  and a_11 (w_11, sel11, data11);
  and a_12 (w_12, sel12, data12);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11, w_12);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux17(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, sel13,
     data13, sel14, data14, sel15, data15, sel16, data16, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12, sel13,
       data13, sel14, data14, sel15, data15, sel16, data16;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12, sel13, data13,
       sel14, data14, sel15, data15, sel16, data16;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or sel9 or sel10 or sel11 or sel12 or sel13 or sel14 or
         sel15 or sel16 or data0 or data1 or data2 or data3 or data4 or
         data5 or data6 or data7 or data8 or data9 or data10 or data11
         or data12 or data13 or data14 or data15 or data16) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
           sel9, sel10, sel11, sel12, sel13, sel14, sel15, sel16})
       17'b10000000000000000: z = data0;
       17'b01000000000000000: z = data1;
       17'b00100000000000000: z = data2;
       17'b00010000000000000: z = data3;
       17'b00001000000000000: z = data4;
       17'b00000100000000000: z = data5;
       17'b00000010000000000: z = data6;
       17'b00000001000000000: z = data7;
       17'b00000000100000000: z = data8;
       17'b00000000010000000: z = data9;
       17'b00000000001000000: z = data10;
       17'b00000000000100000: z = data11;
       17'b00000000000010000: z = data12;
       17'b00000000000001000: z = data13;
       17'b00000000000000100: z = data14;
       17'b00000000000000010: z = data15;
       17'b00000000000000001: z = data16;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux17(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, sel13,
     data13, sel14, data14, sel15, data15, sel16, data16, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12, sel13,
       data13, sel14, data14, sel15, data15, sel16, data16;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12, sel13, data13,
       sel14, data14, sel15, data15, sel16, data16;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8, w_9, w_10, w_11, w_12, w_13, w_14, w_15;
  wire w_16;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  and a_9 (w_9, sel9, data9);
  and a_10 (w_10, sel10, data10);
  and a_11 (w_11, sel11, data11);
  and a_12 (w_12, sel12, data12);
  and a_13 (w_13, sel13, data13);
  and a_14 (w_14, sel14, data14);
  and a_15 (w_15, sel15, data15);
  and a_16 (w_16, sel16, data16);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11, w_12, w_13, w_14, w_15, w_16);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX // captures one-hot property of select inputs
module CDN_mux14(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, sel13,
     data13, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12, sel13,
       data13;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12, sel13, data13;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or sel5 or sel6 or sel7 or
         sel8 or sel9 or sel10 or sel11 or sel12 or sel13 or data0 or
         data1 or data2 or data3 or data4 or data5 or data6 or data7 or
         data8 or data9 or data10 or data11 or data12 or data13) 
      case ({sel0, sel1, sel2, sel3, sel4, sel5, sel6, sel7, sel8,
           sel9, sel10, sel11, sel12, sel13})
       14'b10000000000000: z = data0;
       14'b01000000000000: z = data1;
       14'b00100000000000: z = data2;
       14'b00010000000000: z = data3;
       14'b00001000000000: z = data4;
       14'b00000100000000: z = data5;
       14'b00000010000000: z = data6;
       14'b00000001000000: z = data7;
       14'b00000000100000: z = data8;
       14'b00000000010000: z = data9;
       14'b00000000001000: z = data10;
       14'b00000000000100: z = data11;
       14'b00000000000010: z = data12;
       14'b00000000000001: z = data13;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_mux14(sel0, data0, sel1, data1, sel2, data2, sel3, data3,
     sel4, data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8,
     sel9, data9, sel10, data10, sel11, data11, sel12, data12, sel13,
     data13, z);
  input sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4,
       data4, sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9,
       data9, sel10, data10, sel11, data11, sel12, data12, sel13,
       data13;
  output z;
  wire sel0, data0, sel1, data1, sel2, data2, sel3, data3, sel4, data4,
       sel5, data5, sel6, data6, sel7, data7, sel8, data8, sel9, data9,
       sel10, data10, sel11, data11, sel12, data12, sel13, data13;
  wire z;
  wire w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7;
  wire w_8, w_9, w_10, w_11, w_12, w_13;
  and a_0 (w_0, sel0, data0);
  and a_1 (w_1, sel1, data1);
  and a_2 (w_2, sel2, data2);
  and a_3 (w_3, sel3, data3);
  and a_4 (w_4, sel4, data4);
  and a_5 (w_5, sel5, data5);
  and a_6 (w_6, sel6, data6);
  and a_7 (w_7, sel7, data7);
  and a_8 (w_8, sel8, data8);
  and a_9 (w_9, sel9, data9);
  and a_10 (w_10, sel10, data10);
  and a_11 (w_11, sel11, data11);
  and a_12 (w_12, sel12, data12);
  and a_13 (w_13, sel13, data13);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11, w_12, w_13);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux2(sel0, data0, data1, z);
  input sel0, data0, data1;
  output z;
  wire sel0, data0, data1;
  reg  z;
  always 
    @(sel0 or data0 or data1) 
      case ({sel0})
       1'b0: z = data0;
       1'b1: z = data1;
      endcase
endmodule
`else
module CDN_bmux2(sel0, data0, data1, z);
  input sel0, data0, data1;
  output z;
  wire sel0, data0, data1;
  wire z;
  wire inv_sel0, w_0, w_1;
  not i_0 (inv_sel0, sel0);
  and a_0 (w_0, inv_sel0, data0);
  and a_1 (w_1, sel0, data1);
  or org (z, w_0, w_1);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux9(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or data0 or data1 or data2 or data3
         or data4 or data5 or data6 or data7 or data8) 
      case ({sel0, sel1, sel2, sel3})
       4'b0000: z = data0;
       4'b1000: z = data1;
       4'b0100: z = data2;
       4'b1100: z = data3;
       4'b0010: z = data4;
       4'b1010: z = data5;
       4'b0110: z = data6;
       4'b1110: z = data7;
       4'b0001: z = data8;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_bmux9(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8;
  wire z;
  wire inv_sel0, inv_sel1, inv_sel2, inv_sel3, w_0, w_1, w_2, w_3;
  wire w_4, w_5, w_6, w_7, w_8;
  not i_0 (inv_sel0, sel0);
  not i_1 (inv_sel1, sel1);
  not i_2 (inv_sel2, sel2);
  not i_3 (inv_sel3, sel3);
  and a_0 (w_0, inv_sel3, inv_sel2, inv_sel1, inv_sel0, data0);
  and a_1 (w_1, inv_sel3, inv_sel2, inv_sel1, sel0, data1);
  and a_2 (w_2, inv_sel3, inv_sel2, sel1, inv_sel0, data2);
  and a_3 (w_3, inv_sel3, inv_sel2, sel1, sel0, data3);
  and a_4 (w_4, inv_sel3, sel2, inv_sel1, inv_sel0, data4);
  and a_5 (w_5, inv_sel3, sel2, inv_sel1, sel0, data5);
  and a_6 (w_6, inv_sel3, sel2, sel1, inv_sel0, data6);
  and a_7 (w_7, inv_sel3, sel2, sel1, sel0, data7);
  and a_8 (w_8, sel3, inv_sel2, inv_sel1, inv_sel0, data8);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux8(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or data0 or data1 or data2 or data3 or data4
         or data5 or data6 or data7) 
      case ({sel0, sel1, sel2})
       3'b000: z = data0;
       3'b100: z = data1;
       3'b010: z = data2;
       3'b110: z = data3;
       3'b001: z = data4;
       3'b101: z = data5;
       3'b011: z = data6;
       3'b111: z = data7;
      endcase
endmodule
`else
module CDN_bmux8(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7;
  wire z;
  wire inv_sel0, inv_sel1, inv_sel2, w_0, w_1, w_2, w_3, w_4;
  wire w_5, w_6, w_7;
  not i_0 (inv_sel0, sel0);
  not i_1 (inv_sel1, sel1);
  not i_2 (inv_sel2, sel2);
  and a_0 (w_0, inv_sel2, inv_sel1, inv_sel0, data0);
  and a_1 (w_1, inv_sel2, inv_sel1, sel0, data1);
  and a_2 (w_2, inv_sel2, sel1, inv_sel0, data2);
  and a_3 (w_3, inv_sel2, sel1, sel0, data3);
  and a_4 (w_4, sel2, inv_sel1, inv_sel0, data4);
  and a_5 (w_5, sel2, inv_sel1, sel0, data5);
  and a_6 (w_6, sel2, sel1, inv_sel0, data6);
  and a_7 (w_7, sel2, sel1, sel0, data7);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux16(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, data9, data10, data11, data12,
     data13, data14, data15, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or data0 or data1 or data2 or data3
         or data4 or data5 or data6 or data7 or data8 or data9 or
         data10 or data11 or data12 or data13 or data14 or data15) 
      case ({sel0, sel1, sel2, sel3})
       4'b0000: z = data0;
       4'b1000: z = data1;
       4'b0100: z = data2;
       4'b1100: z = data3;
       4'b0010: z = data4;
       4'b1010: z = data5;
       4'b0110: z = data6;
       4'b1110: z = data7;
       4'b0001: z = data8;
       4'b1001: z = data9;
       4'b0101: z = data10;
       4'b1101: z = data11;
       4'b0011: z = data12;
       4'b1011: z = data13;
       4'b0111: z = data14;
       4'b1111: z = data15;
      endcase
endmodule
`else
module CDN_bmux16(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, data9, data10, data11, data12,
     data13, data14, data15, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15;
  wire z;
  wire inv_sel0, inv_sel1, inv_sel2, inv_sel3, w_0, w_1, w_2, w_3;
  wire w_4, w_5, w_6, w_7, w_8, w_9, w_10, w_11;
  wire w_12, w_13, w_14, w_15;
  not i_0 (inv_sel0, sel0);
  not i_1 (inv_sel1, sel1);
  not i_2 (inv_sel2, sel2);
  not i_3 (inv_sel3, sel3);
  and a_0 (w_0, inv_sel3, inv_sel2, inv_sel1, inv_sel0, data0);
  and a_1 (w_1, inv_sel3, inv_sel2, inv_sel1, sel0, data1);
  and a_2 (w_2, inv_sel3, inv_sel2, sel1, inv_sel0, data2);
  and a_3 (w_3, inv_sel3, inv_sel2, sel1, sel0, data3);
  and a_4 (w_4, inv_sel3, sel2, inv_sel1, inv_sel0, data4);
  and a_5 (w_5, inv_sel3, sel2, inv_sel1, sel0, data5);
  and a_6 (w_6, inv_sel3, sel2, sel1, inv_sel0, data6);
  and a_7 (w_7, inv_sel3, sel2, sel1, sel0, data7);
  and a_8 (w_8, sel3, inv_sel2, inv_sel1, inv_sel0, data8);
  and a_9 (w_9, sel3, inv_sel2, inv_sel1, sel0, data9);
  and a_10 (w_10, sel3, inv_sel2, sel1, inv_sel0, data10);
  and a_11 (w_11, sel3, inv_sel2, sel1, sel0, data11);
  and a_12 (w_12, sel3, sel2, inv_sel1, inv_sel0, data12);
  and a_13 (w_13, sel3, sel2, inv_sel1, sel0, data13);
  and a_14 (w_14, sel3, sel2, sel1, inv_sel0, data14);
  and a_15 (w_15, sel3, sel2, sel1, sel0, data15);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11, w_12, w_13, w_14, w_15);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux7(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or data0 or data1 or data2 or data3 or data4
         or data5 or data6) 
      case ({sel0, sel1, sel2})
       3'b000: z = data0;
       3'b100: z = data1;
       3'b010: z = data2;
       3'b110: z = data3;
       3'b001: z = data4;
       3'b101: z = data5;
       3'b011: z = data6;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_bmux7(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6;
  wire z;
  wire inv_sel0, inv_sel1, inv_sel2, w_0, w_1, w_2, w_3, w_4;
  wire w_5, w_6;
  not i_0 (inv_sel0, sel0);
  not i_1 (inv_sel1, sel1);
  not i_2 (inv_sel2, sel2);
  and a_0 (w_0, inv_sel2, inv_sel1, inv_sel0, data0);
  and a_1 (w_1, inv_sel2, inv_sel1, sel0, data1);
  and a_2 (w_2, inv_sel2, sel1, inv_sel0, data2);
  and a_3 (w_3, inv_sel2, sel1, sel0, data3);
  and a_4 (w_4, sel2, inv_sel1, inv_sel0, data4);
  and a_5 (w_5, sel2, inv_sel1, sel0, data5);
  and a_6 (w_6, sel2, sel1, inv_sel0, data6);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux4(sel0, data0, data1, sel1, data2, data3, z);
  input sel0, data0, data1, sel1, data2, data3;
  output z;
  wire sel0, data0, data1, sel1, data2, data3;
  reg  z;
  always 
    @(sel0 or sel1 or data0 or data1 or data2 or data3) 
      case ({sel0, sel1})
       2'b00: z = data0;
       2'b10: z = data1;
       2'b01: z = data2;
       2'b11: z = data3;
      endcase
endmodule
`else
module CDN_bmux4(sel0, data0, data1, sel1, data2, data3, z);
  input sel0, data0, data1, sel1, data2, data3;
  output z;
  wire sel0, data0, data1, sel1, data2, data3;
  wire z;
  wire inv_sel0, inv_sel1, w_0, w_1, w_2, w_3;
  not i_0 (inv_sel0, sel0);
  not i_1 (inv_sel1, sel1);
  and a_0 (w_0, inv_sel1, inv_sel0, data0);
  and a_1 (w_1, inv_sel1, sel0, data1);
  and a_2 (w_2, sel1, inv_sel0, data2);
  and a_3 (w_3, sel1, sel0, data3);
  or org (z, w_0, w_1, w_2, w_3);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux31(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, data9, data10, data11, data12,
     data13, data14, data15, sel4, data16, data17, data18, data19,
     data20, data21, data22, data23, data24, data25, data26, data27,
     data28, data29, data30, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17, data18, data19,
       data20, data21, data22, data23, data24, data25, data26, data27,
       data28, data29, data30;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17, data18, data19,
       data20, data21, data22, data23, data24, data25, data26, data27,
       data28, data29, data30;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or data0 or data1 or data2
         or data3 or data4 or data5 or data6 or data7 or data8 or data9
         or data10 or data11 or data12 or data13 or data14 or data15 or
         data16 or data17 or data18 or data19 or data20 or data21 or
         data22 or data23 or data24 or data25 or data26 or data27 or
         data28 or data29 or data30) 
      case ({sel0, sel1, sel2, sel3, sel4})
       5'b00000: z = data0;
       5'b10000: z = data1;
       5'b01000: z = data2;
       5'b11000: z = data3;
       5'b00100: z = data4;
       5'b10100: z = data5;
       5'b01100: z = data6;
       5'b11100: z = data7;
       5'b00010: z = data8;
       5'b10010: z = data9;
       5'b01010: z = data10;
       5'b11010: z = data11;
       5'b00110: z = data12;
       5'b10110: z = data13;
       5'b01110: z = data14;
       5'b11110: z = data15;
       5'b00001: z = data16;
       5'b10001: z = data17;
       5'b01001: z = data18;
       5'b11001: z = data19;
       5'b00101: z = data20;
       5'b10101: z = data21;
       5'b01101: z = data22;
       5'b11101: z = data23;
       5'b00011: z = data24;
       5'b10011: z = data25;
       5'b01011: z = data26;
       5'b11011: z = data27;
       5'b00111: z = data28;
       5'b10111: z = data29;
       5'b01111: z = data30;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_bmux31(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, data9, data10, data11, data12,
     data13, data14, data15, sel4, data16, data17, data18, data19,
     data20, data21, data22, data23, data24, data25, data26, data27,
     data28, data29, data30, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17, data18, data19,
       data20, data21, data22, data23, data24, data25, data26, data27,
       data28, data29, data30;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17, data18, data19,
       data20, data21, data22, data23, data24, data25, data26, data27,
       data28, data29, data30;
  wire z;
  wire inv_sel0, inv_sel1, inv_sel2, inv_sel3, inv_sel4, w_0, w_1, w_2;
  wire w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10;
  wire w_11, w_12, w_13, w_14, w_15, w_16, w_17, w_18;
  wire w_19, w_20, w_21, w_22, w_23, w_24, w_25, w_26;
  wire w_27, w_28, w_29, w_30;
  not i_0 (inv_sel0, sel0);
  not i_1 (inv_sel1, sel1);
  not i_2 (inv_sel2, sel2);
  not i_3 (inv_sel3, sel3);
  not i_4 (inv_sel4, sel4);
  and a_0 (w_0, inv_sel4, inv_sel3, inv_sel2, inv_sel1, inv_sel0,
       data0);
  and a_1 (w_1, inv_sel4, inv_sel3, inv_sel2, inv_sel1, sel0, data1);
  and a_2 (w_2, inv_sel4, inv_sel3, inv_sel2, sel1, inv_sel0, data2);
  and a_3 (w_3, inv_sel4, inv_sel3, inv_sel2, sel1, sel0, data3);
  and a_4 (w_4, inv_sel4, inv_sel3, sel2, inv_sel1, inv_sel0, data4);
  and a_5 (w_5, inv_sel4, inv_sel3, sel2, inv_sel1, sel0, data5);
  and a_6 (w_6, inv_sel4, inv_sel3, sel2, sel1, inv_sel0, data6);
  and a_7 (w_7, inv_sel4, inv_sel3, sel2, sel1, sel0, data7);
  and a_8 (w_8, inv_sel4, sel3, inv_sel2, inv_sel1, inv_sel0, data8);
  and a_9 (w_9, inv_sel4, sel3, inv_sel2, inv_sel1, sel0, data9);
  and a_10 (w_10, inv_sel4, sel3, inv_sel2, sel1, inv_sel0, data10);
  and a_11 (w_11, inv_sel4, sel3, inv_sel2, sel1, sel0, data11);
  and a_12 (w_12, inv_sel4, sel3, sel2, inv_sel1, inv_sel0, data12);
  and a_13 (w_13, inv_sel4, sel3, sel2, inv_sel1, sel0, data13);
  and a_14 (w_14, inv_sel4, sel3, sel2, sel1, inv_sel0, data14);
  and a_15 (w_15, inv_sel4, sel3, sel2, sel1, sel0, data15);
  and a_16 (w_16, sel4, inv_sel3, inv_sel2, inv_sel1, inv_sel0, data16);
  and a_17 (w_17, sel4, inv_sel3, inv_sel2, inv_sel1, sel0, data17);
  and a_18 (w_18, sel4, inv_sel3, inv_sel2, sel1, inv_sel0, data18);
  and a_19 (w_19, sel4, inv_sel3, inv_sel2, sel1, sel0, data19);
  and a_20 (w_20, sel4, inv_sel3, sel2, inv_sel1, inv_sel0, data20);
  and a_21 (w_21, sel4, inv_sel3, sel2, inv_sel1, sel0, data21);
  and a_22 (w_22, sel4, inv_sel3, sel2, sel1, inv_sel0, data22);
  and a_23 (w_23, sel4, inv_sel3, sel2, sel1, sel0, data23);
  and a_24 (w_24, sel4, sel3, inv_sel2, inv_sel1, inv_sel0, data24);
  and a_25 (w_25, sel4, sel3, inv_sel2, inv_sel1, sel0, data25);
  and a_26 (w_26, sel4, sel3, inv_sel2, sel1, inv_sel0, data26);
  and a_27 (w_27, sel4, sel3, inv_sel2, sel1, sel0, data27);
  and a_28 (w_28, sel4, sel3, sel2, inv_sel1, inv_sel0, data28);
  and a_29 (w_29, sel4, sel3, sel2, inv_sel1, sel0, data29);
  and a_30 (w_30, sel4, sel3, sel2, sel1, inv_sel0, data30);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11, w_12, w_13, w_14, w_15, w_16, w_17, w_18, w_19, w_20,
       w_21, w_22, w_23, w_24, w_25, w_26, w_27, w_28, w_29, w_30);
endmodule
`endif // ONE_HOT_MUX
`endif
`ifdef RC_CDN_GENERIC_GATE
`else
`ifdef ONE_HOT_MUX
module CDN_bmux18(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, data9, data10, data11, data12,
     data13, data14, data15, sel4, data16, data17, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17;
  reg  z;
  always 
    @(sel0 or sel1 or sel2 or sel3 or sel4 or data0 or data1 or data2
         or data3 or data4 or data5 or data6 or data7 or data8 or data9
         or data10 or data11 or data12 or data13 or data14 or data15 or
         data16 or data17) 
      case ({sel0, sel1, sel2, sel3, sel4})
       5'b00000: z = data0;
       5'b10000: z = data1;
       5'b01000: z = data2;
       5'b11000: z = data3;
       5'b00100: z = data4;
       5'b10100: z = data5;
       5'b01100: z = data6;
       5'b11100: z = data7;
       5'b00010: z = data8;
       5'b10010: z = data9;
       5'b01010: z = data10;
       5'b11010: z = data11;
       5'b00110: z = data12;
       5'b10110: z = data13;
       5'b01110: z = data14;
       5'b11110: z = data15;
       5'b00001: z = data16;
       5'b10001: z = data17;
       default: z = 1'bX;
      endcase
endmodule
`else
module CDN_bmux18(sel0, data0, data1, sel1, data2, data3, sel2, data4,
     data5, data6, data7, sel3, data8, data9, data10, data11, data12,
     data13, data14, data15, sel4, data16, data17, z);
  input sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17;
  output z;
  wire sel0, data0, data1, sel1, data2, data3, sel2, data4, data5,
       data6, data7, sel3, data8, data9, data10, data11, data12,
       data13, data14, data15, sel4, data16, data17;
  wire z;
  wire inv_sel0, inv_sel1, inv_sel2, inv_sel3, inv_sel4, w_0, w_1, w_2;
  wire w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10;
  wire w_11, w_12, w_13, w_14, w_15, w_16, w_17;
  not i_0 (inv_sel0, sel0);
  not i_1 (inv_sel1, sel1);
  not i_2 (inv_sel2, sel2);
  not i_3 (inv_sel3, sel3);
  not i_4 (inv_sel4, sel4);
  and a_0 (w_0, inv_sel4, inv_sel3, inv_sel2, inv_sel1, inv_sel0,
       data0);
  and a_1 (w_1, inv_sel4, inv_sel3, inv_sel2, inv_sel1, sel0, data1);
  and a_2 (w_2, inv_sel4, inv_sel3, inv_sel2, sel1, inv_sel0, data2);
  and a_3 (w_3, inv_sel4, inv_sel3, inv_sel2, sel1, sel0, data3);
  and a_4 (w_4, inv_sel4, inv_sel3, sel2, inv_sel1, inv_sel0, data4);
  and a_5 (w_5, inv_sel4, inv_sel3, sel2, inv_sel1, sel0, data5);
  and a_6 (w_6, inv_sel4, inv_sel3, sel2, sel1, inv_sel0, data6);
  and a_7 (w_7, inv_sel4, inv_sel3, sel2, sel1, sel0, data7);
  and a_8 (w_8, inv_sel4, sel3, inv_sel2, inv_sel1, inv_sel0, data8);
  and a_9 (w_9, inv_sel4, sel3, inv_sel2, inv_sel1, sel0, data9);
  and a_10 (w_10, inv_sel4, sel3, inv_sel2, sel1, inv_sel0, data10);
  and a_11 (w_11, inv_sel4, sel3, inv_sel2, sel1, sel0, data11);
  and a_12 (w_12, inv_sel4, sel3, sel2, inv_sel1, inv_sel0, data12);
  and a_13 (w_13, inv_sel4, sel3, sel2, inv_sel1, sel0, data13);
  and a_14 (w_14, inv_sel4, sel3, sel2, sel1, inv_sel0, data14);
  and a_15 (w_15, inv_sel4, sel3, sel2, sel1, sel0, data15);
  and a_16 (w_16, sel4, inv_sel3, inv_sel2, inv_sel1, inv_sel0, data16);
  and a_17 (w_17, sel4, inv_sel3, inv_sel2, inv_sel1, sel0, data17);
  or org (z, w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10,
       w_11, w_12, w_13, w_14, w_15, w_16, w_17);
endmodule
`endif // ONE_HOT_MUX
`endif
