//
// FX68K
//
// M68K cycle accurate, fully synchronous
// Copyright 2018 by Jorge Cwik
//
module uRom( input clk, input [10-1:0] microAddr, output reg [17-1:0] microOutput);

  always @( posedge clk)
  begin
    case (microAddr)
      10'h  0 : microOutput = 17'b10010000101100000;
      10'h  1 : microOutput = 17'b10000100000000000;
      10'h  2 : microOutput = 17'b00101001011010000;
      10'h  3 : microOutput = 17'b00111110011000000;
      10'h  4 : microOutput = 17'b01000000000001100;
      10'h  5 : microOutput = 17'b01000000000001100;
      10'h  6 : microOutput = 17'b01000010010000000;
      10'h  7 : microOutput = 17'b10001100011100000;
      10'h  8 : microOutput = 17'b01000100010000000;
      10'h  9 : microOutput = 17'b10000000010000000;
      10'h  a : microOutput = 17'b10000000010000000;
      10'h  b : microOutput = 17'b01000100010000000;
      10'h  c : microOutput = 17'b00001010010000000;
      10'h  d : microOutput = 17'b10000000100000000;
      10'h  e : microOutput = 17'b10000000100000000;
      10'h  f : microOutput = 17'b01101001100000000;
      10'h 10 : microOutput = 17'b00000000000000000;
      10'h 11 : microOutput = 17'b00000000000000000;
      10'h 12 : microOutput = 17'b00000000000000000;
      10'h 13 : microOutput = 17'b00000000000000000;
      10'h 14 : microOutput = 17'b00000000000000000;
      10'h 15 : microOutput = 17'b00000000000000000;
      10'h 16 : microOutput = 17'b00000000000000000;
      10'h 17 : microOutput = 17'b00000000000000000;
      10'h 18 : microOutput = 17'b00000000000000000;
      10'h 19 : microOutput = 17'b00000000000000000;
      10'h 1a : microOutput = 17'b00000000000000000;
      10'h 1b : microOutput = 17'b00000000000000000;
      10'h 1c : microOutput = 17'b00000000000000000;
      10'h 1d : microOutput = 17'b00000000000000000;
      10'h 1e : microOutput = 17'b00000000000000000;
      10'h 1f : microOutput = 17'b00000000000000000;
      10'h 20 : microOutput = 17'b00000000000000100;
      10'h 21 : microOutput = 17'b00001010110000000;
      10'h 22 : microOutput = 17'b00111000001100000;
      10'h 23 : microOutput = 17'b00100101001001010;
      10'h 24 : microOutput = 17'b00000000000001100;
      10'h 25 : microOutput = 17'b10110000110100001;
      10'h 26 : microOutput = 17'b00000000000001100;
      10'h 27 : microOutput = 17'b00001110100000000;
      10'h 28 : microOutput = 17'b00110100101000000;
      10'h 29 : microOutput = 17'b00100011010100000;
      10'h 2a : microOutput = 17'b00000010010000000;
      10'h 2b : microOutput = 17'b10000110000000010;
      10'h 2c : microOutput = 17'b00111110110000000;
      10'h 2d : microOutput = 17'b00000100011100000;
      10'h 2e : microOutput = 17'b00101111010100000;
      10'h 2f : microOutput = 17'b10010011100000010;
      10'h 30 : microOutput = 17'b00000000000000000;
      10'h 31 : microOutput = 17'b00000000000000000;
      10'h 32 : microOutput = 17'b00000000000000000;
      10'h 33 : microOutput = 17'b00000000000000000;
      10'h 34 : microOutput = 17'b00000000000000000;
      10'h 35 : microOutput = 17'b00000000000000000;
      10'h 36 : microOutput = 17'b00000000000000000;
      10'h 37 : microOutput = 17'b00000000000000000;
      10'h 38 : microOutput = 17'b00000000000000000;
      10'h 39 : microOutput = 17'b00000000000000000;
      10'h 3a : microOutput = 17'b00000000000000000;
      10'h 3b : microOutput = 17'b00000000000000000;
      10'h 3c : microOutput = 17'b00000000000000000;
      10'h 3d : microOutput = 17'b00000000000000000;
      10'h 3e : microOutput = 17'b00000000000000000;
      10'h 3f : microOutput = 17'b00000000000000000;
      10'h 40 : microOutput = 17'b10011101000000000;
      10'h 41 : microOutput = 17'b00000100110010110;
      10'h 42 : microOutput = 17'b00101001010000000;
      10'h 43 : microOutput = 17'b10110000110100001;
      10'h 44 : microOutput = 17'b00000000000000100;
      10'h 45 : microOutput = 17'b00111110000100000;
      10'h 46 : microOutput = 17'b10010111010100000;
      10'h 47 : microOutput = 17'b01000110000100000;
      10'h 48 : microOutput = 17'b01010111100000000;
      10'h 49 : microOutput = 17'b10001010010011010;
      10'h 4a : microOutput = 17'b01000110010100001;
      10'h 4b : microOutput = 17'b00000110010111010;
      10'h 4c : microOutput = 17'b01001100010100000;
      10'h 4d : microOutput = 17'b10001010010010111;
      10'h 4e : microOutput = 17'b01000000000100001;
      10'h 4f : microOutput = 17'b00110100111000000;
      10'h 50 : microOutput = 17'b00000000000000000;
      10'h 51 : microOutput = 17'b00000000000000000;
      10'h 52 : microOutput = 17'b00000000000000000;
      10'h 53 : microOutput = 17'b00000000000000000;
      10'h 54 : microOutput = 17'b00000000000000000;
      10'h 55 : microOutput = 17'b00000000000000000;
      10'h 56 : microOutput = 17'b00000000000000000;
      10'h 57 : microOutput = 17'b00000000000000000;
      10'h 58 : microOutput = 17'b00000000000000000;
      10'h 59 : microOutput = 17'b00000000000000000;
      10'h 5a : microOutput = 17'b00000000000000000;
      10'h 5b : microOutput = 17'b00000000000000000;
      10'h 5c : microOutput = 17'b00000000000000000;
      10'h 5d : microOutput = 17'b00000000000000000;
      10'h 5e : microOutput = 17'b00000000000000000;
      10'h 5f : microOutput = 17'b00000000000000000;
      10'h 60 : microOutput = 17'b00000010001100000;
      10'h 61 : microOutput = 17'b01001010000100001;
      10'h 62 : microOutput = 17'b10110100111000000;
      10'h 63 : microOutput = 17'b00011011010100000;
      10'h 64 : microOutput = 17'b10000000000000100;
      10'h 65 : microOutput = 17'b10110100111000000;
      10'h 66 : microOutput = 17'b00000000000000100;
      10'h 67 : microOutput = 17'b00001000001000000;
      10'h 68 : microOutput = 17'b00000100011100110;
      10'h 69 : microOutput = 17'b10001110010100001;
      10'h 6a : microOutput = 17'b00000000011110010;
      10'h 6b : microOutput = 17'b01001000011000000;
      10'h 6c : microOutput = 17'b00001000010100110;
      10'h 6d : microOutput = 17'b10001010000110111;
      10'h 6e : microOutput = 17'b00000000111110010;
      10'h 6f : microOutput = 17'b01001000111000000;
      10'h 70 : microOutput = 17'b00000000000000000;
      10'h 71 : microOutput = 17'b00000000000000000;
      10'h 72 : microOutput = 17'b00000000000000000;
      10'h 73 : microOutput = 17'b00000000000000000;
      10'h 74 : microOutput = 17'b00000000000000000;
      10'h 75 : microOutput = 17'b00000000000000000;
      10'h 76 : microOutput = 17'b00000000000000000;
      10'h 77 : microOutput = 17'b00000000000000000;
      10'h 78 : microOutput = 17'b00000000000000000;
      10'h 79 : microOutput = 17'b00000000000000000;
      10'h 7a : microOutput = 17'b00000000000000000;
      10'h 7b : microOutput = 17'b00000000000000000;
      10'h 7c : microOutput = 17'b00000000000000000;
      10'h 7d : microOutput = 17'b00000000000000000;
      10'h 7e : microOutput = 17'b00000000000000000;
      10'h 7f : microOutput = 17'b00000000000000000;
      10'h 80 : microOutput = 17'b10101001000000001;
      10'h 81 : microOutput = 17'b10001000001000001;
      10'h 82 : microOutput = 17'b01000000000000100;
      10'h 83 : microOutput = 17'b01001100001111010;
      10'h 84 : microOutput = 17'b00000110001000000;
      10'h 85 : microOutput = 17'b00010110001100000;
      10'h 86 : microOutput = 17'b00011010000000000;
      10'h 87 : microOutput = 17'b10110000110100001;
      10'h 88 : microOutput = 17'b01111000001100000;
      10'h 89 : microOutput = 17'b00011000000000000;
      10'h 8a : microOutput = 17'b00000100100100001;
      10'h 8b : microOutput = 17'b00000000000000100;
      10'h 8c : microOutput = 17'b00000000101100000;
      10'h 8d : microOutput = 17'b00000000000000100;
      10'h 8e : microOutput = 17'b00010001010100000;
      10'h 8f : microOutput = 17'b10010111000100001;
      10'h 90 : microOutput = 17'b00000000000000000;
      10'h 91 : microOutput = 17'b00000000000000000;
      10'h 92 : microOutput = 17'b00000000000000000;
      10'h 93 : microOutput = 17'b00000000000000000;
      10'h 94 : microOutput = 17'b00000000000000000;
      10'h 95 : microOutput = 17'b00000000000000000;
      10'h 96 : microOutput = 17'b00000000000000000;
      10'h 97 : microOutput = 17'b00000000000000000;
      10'h 98 : microOutput = 17'b00000000000000000;
      10'h 99 : microOutput = 17'b00000000000000000;
      10'h 9a : microOutput = 17'b00000000000000000;
      10'h 9b : microOutput = 17'b00000000000000000;
      10'h 9c : microOutput = 17'b00000000000000000;
      10'h 9d : microOutput = 17'b00000000000000000;
      10'h 9e : microOutput = 17'b00000000000000000;
      10'h 9f : microOutput = 17'b00000000000000000;
      10'h a0 : microOutput = 17'b00000010001100000;
      10'h a1 : microOutput = 17'b00000000000000100;
      10'h a2 : microOutput = 17'b01111000011100000;
      10'h a3 : microOutput = 17'b00011011010100000;
      10'h a4 : microOutput = 17'b00101101000000000;
      10'h a5 : microOutput = 17'b01000110010111010;
      10'h a6 : microOutput = 17'b00101101000000000;
      10'h a7 : microOutput = 17'b10001010101100000;
      10'h a8 : microOutput = 17'b01010110001100000;
      10'h a9 : microOutput = 17'b00011000110000000;
      10'h aa : microOutput = 17'b01010110001100000;
      10'h ab : microOutput = 17'b10001110011100001;
      10'h ac : microOutput = 17'b00000100101100000;
      10'h ad : microOutput = 17'b01000110010111010;
      10'h ae : microOutput = 17'b00000100101100000;
      10'h af : microOutput = 17'b10001010111100000;
      10'h b0 : microOutput = 17'b00000000000000000;
      10'h b1 : microOutput = 17'b00000000000000000;
      10'h b2 : microOutput = 17'b00000000000000000;
      10'h b3 : microOutput = 17'b00000000000000000;
      10'h b4 : microOutput = 17'b00000000000000000;
      10'h b5 : microOutput = 17'b00000000000000000;
      10'h b6 : microOutput = 17'b00000000000000000;
      10'h b7 : microOutput = 17'b00000000000000000;
      10'h b8 : microOutput = 17'b00000000000000000;
      10'h b9 : microOutput = 17'b00000000000000000;
      10'h ba : microOutput = 17'b00000000000000000;
      10'h bb : microOutput = 17'b00000000000000000;
      10'h bc : microOutput = 17'b00000000000000000;
      10'h bd : microOutput = 17'b00000000000000000;
      10'h be : microOutput = 17'b00000000000000000;
      10'h bf : microOutput = 17'b00000000000000000;
      10'h c0 : microOutput = 17'b10101001000000001;
      10'h c1 : microOutput = 17'b00001000101010110;
      10'h c2 : microOutput = 17'b00011111010100000;
      10'h c3 : microOutput = 17'b01101101110000000;
      10'h c4 : microOutput = 17'b00000000000000100;
      10'h c5 : microOutput = 17'b10111110000100000;
      10'h c6 : microOutput = 17'b00000100011100000;
      10'h c7 : microOutput = 17'b10001100101000001;
      10'h c8 : microOutput = 17'b00000110001000000;
      10'h c9 : microOutput = 17'b00001110000010010;
      10'h ca : microOutput = 17'b00100101000010110;
      10'h cb : microOutput = 17'b00101101000100000;
      10'h cc : microOutput = 17'b00000000011100000;
      10'h cd : microOutput = 17'b00001000111100000;
      10'h ce : microOutput = 17'b00100101000011010;
      10'h cf : microOutput = 17'b00110100111000000;
      10'h d0 : microOutput = 17'b00000000000000000;
      10'h d1 : microOutput = 17'b00000000000000000;
      10'h d2 : microOutput = 17'b00000000000000000;
      10'h d3 : microOutput = 17'b00000000000000000;
      10'h d4 : microOutput = 17'b00000000000000000;
      10'h d5 : microOutput = 17'b00000000000000000;
      10'h d6 : microOutput = 17'b00000000000000000;
      10'h d7 : microOutput = 17'b00000000000000000;
      10'h d8 : microOutput = 17'b00000000000000000;
      10'h d9 : microOutput = 17'b00000000000000000;
      10'h da : microOutput = 17'b00000000000000000;
      10'h db : microOutput = 17'b00000000000000000;
      10'h dc : microOutput = 17'b00000000000000000;
      10'h dd : microOutput = 17'b00000000000000000;
      10'h de : microOutput = 17'b00000000000000000;
      10'h df : microOutput = 17'b00000000000000000;
      10'h e0 : microOutput = 17'b00000010000100010;
      10'h e1 : microOutput = 17'b00001010110000000;
      10'h e2 : microOutput = 17'b00000000000000100;
      10'h e3 : microOutput = 17'b00101101010000000;
      10'h e4 : microOutput = 17'b01010001010000000;
      10'h e5 : microOutput = 17'b01000110111000000;
      10'h e6 : microOutput = 17'b00000000000000100;
      10'h e7 : microOutput = 17'b00000000010110010;
      10'h e8 : microOutput = 17'b00110100101000000;
      10'h e9 : microOutput = 17'b00100011010100000;
      10'h ea : microOutput = 17'b10000000000001000;
      10'h eb : microOutput = 17'b01101011010000000;
      10'h ec : microOutput = 17'b00111110110000000;
      10'h ed : microOutput = 17'b00000100011100000;
      10'h ee : microOutput = 17'b10010101000000000;
      10'h ef : microOutput = 17'b01111110010100000;
      10'h f0 : microOutput = 17'b00000000000000000;
      10'h f1 : microOutput = 17'b00000000000000000;
      10'h f2 : microOutput = 17'b00000000000000000;
      10'h f3 : microOutput = 17'b00000000000000000;
      10'h f4 : microOutput = 17'b00000000000000000;
      10'h f5 : microOutput = 17'b00000000000000000;
      10'h f6 : microOutput = 17'b00000000000000000;
      10'h f7 : microOutput = 17'b00000000000000000;
      10'h f8 : microOutput = 17'b00000000000000000;
      10'h f9 : microOutput = 17'b00000000000000000;
      10'h fa : microOutput = 17'b00000000000000000;
      10'h fb : microOutput = 17'b00000000000000000;
      10'h fc : microOutput = 17'b00000000000000000;
      10'h fd : microOutput = 17'b00000000000000000;
      10'h fe : microOutput = 17'b00000000000000000;
      10'h ff : microOutput = 17'b00000000000000000;
      10'h100 : microOutput = 17'b10001100101000001;
      10'h101 : microOutput = 17'b10000010100000010;
      10'h102 : microOutput = 17'b01000010101000000;
      10'h103 : microOutput = 17'b00011111100100000;
      10'h104 : microOutput = 17'b10100111100000001;
      10'h105 : microOutput = 17'b10010010110000010;
      10'h106 : microOutput = 17'b01110100111000000;
      10'h107 : microOutput = 17'b00010111010000000;
      10'h108 : microOutput = 17'b10101011100000001;
      10'h109 : microOutput = 17'b10010010100000010;
      10'h10a : microOutput = 17'b01110000100100000;
      10'h10b : microOutput = 17'b00000000100100000;
      10'h10c : microOutput = 17'b10100101100100001;
      10'h10d : microOutput = 17'b10000010110000010;
      10'h10e : microOutput = 17'b01001010101000000;
      10'h10f : microOutput = 17'b00010111000000000;
      10'h110 : microOutput = 17'b00010001000010110;
      10'h111 : microOutput = 17'b01110010100111010;
      10'h112 : microOutput = 17'b10110100010000000;
      10'h113 : microOutput = 17'b00110100111000000;
      10'h114 : microOutput = 17'b01000010010000110;
      10'h115 : microOutput = 17'b01110010110111011;
      10'h116 : microOutput = 17'b01111100000000000;
      10'h117 : microOutput = 17'b00101101000100000;
      10'h118 : microOutput = 17'b00101001001010001;
      10'h119 : microOutput = 17'b01011011111100000;
      10'h11a : microOutput = 17'b01101111011000000;
      10'h11b : microOutput = 17'b00100011100000000;
      10'h11c : microOutput = 17'b00111110000110000;
      10'h11d : microOutput = 17'b00000000000000000;
      10'h11e : microOutput = 17'b10101111011000000;
      10'h11f : microOutput = 17'b00000000000000000;
      10'h120 : microOutput = 17'b00001010100000000;
      10'h121 : microOutput = 17'b10101011100100001;
      10'h122 : microOutput = 17'b01010011000100001;
      10'h123 : microOutput = 17'b10010101010000000;
      10'h124 : microOutput = 17'b00000000110000000;
      10'h125 : microOutput = 17'b10111010000100001;
      10'h126 : microOutput = 17'b01011001010000000;
      10'h127 : microOutput = 17'b10010101000000000;
      10'h128 : microOutput = 17'b00101101101100000;
      10'h129 : microOutput = 17'b10100011100100001;
      10'h12a : microOutput = 17'b01011110100000000;
      10'h12b : microOutput = 17'b01110100011100000;
      10'h12c : microOutput = 17'b00101011111000000;
      10'h12d : microOutput = 17'b10110000110100001;
      10'h12e : microOutput = 17'b01010101010100001;
      10'h12f : microOutput = 17'b00000000000000000;
      10'h130 : microOutput = 17'b00111000100000000;
      10'h131 : microOutput = 17'b01011011000000000;
      10'h132 : microOutput = 17'b00001000100100000;
      10'h133 : microOutput = 17'b10001100101000001;
      10'h134 : microOutput = 17'b00100001100000000;
      10'h135 : microOutput = 17'b01011011010000000;
      10'h136 : microOutput = 17'b00001000110100000;
      10'h137 : microOutput = 17'b10011001110100001;
      10'h138 : microOutput = 17'b00000110010111010;
      10'h139 : microOutput = 17'b01011011100000000;
      10'h13a : microOutput = 17'b00000000110100000;
      10'h13b : microOutput = 17'b10011101010000001;
      10'h13c : microOutput = 17'b00000000000000000;
      10'h13d : microOutput = 17'b00000000000000000;
      10'h13e : microOutput = 17'b00000000000000000;
      10'h13f : microOutput = 17'b00000000000000000;
      10'h140 : microOutput = 17'b00000000000000000;
      10'h141 : microOutput = 17'b00000000000000000;
      10'h142 : microOutput = 17'b00000000000000000;
      10'h143 : microOutput = 17'b00000000000000000;
      10'h144 : microOutput = 17'b00000000000000000;
      10'h145 : microOutput = 17'b00000000000000000;
      10'h146 : microOutput = 17'b00000000000000000;
      10'h147 : microOutput = 17'b00000000000000000;
      10'h148 : microOutput = 17'b00000000000000000;
      10'h149 : microOutput = 17'b00000000000000000;
      10'h14a : microOutput = 17'b00000000000000000;
      10'h14b : microOutput = 17'b00000000000000000;
      10'h14c : microOutput = 17'b00000000000000000;
      10'h14d : microOutput = 17'b00000000000000000;
      10'h14e : microOutput = 17'b00000000000000000;
      10'h14f : microOutput = 17'b00000000000000000;
      10'h150 : microOutput = 17'b10110000110100001;
      10'h151 : microOutput = 17'b00011101000100000;
      10'h152 : microOutput = 17'b00011101000100000;
      10'h153 : microOutput = 17'b00010001000101110;
      10'h154 : microOutput = 17'b01011010110000000;
      10'h155 : microOutput = 17'b01011001010100000;
      10'h156 : microOutput = 17'b10011101010100000;
      10'h157 : microOutput = 17'b00000000000000100;
      10'h158 : microOutput = 17'b10110000110100001;
      10'h159 : microOutput = 17'b00110110000000000;
      10'h15a : microOutput = 17'b10110000011100001;
      10'h15b : microOutput = 17'b10110000011100001;
      10'h15c : microOutput = 17'b10011101000000001;
      10'h15d : microOutput = 17'b01110100111000000;
      10'h15e : microOutput = 17'b00101101100100000;
      10'h15f : microOutput = 17'b10011000100000000;
      10'h160 : microOutput = 17'b00000000000000000;
      10'h161 : microOutput = 17'b00000000000000000;
      10'h162 : microOutput = 17'b00000000000000000;
      10'h163 : microOutput = 17'b00000000000000000;
      10'h164 : microOutput = 17'b00000000000000000;
      10'h165 : microOutput = 17'b00000000000000000;
      10'h166 : microOutput = 17'b00000000000000000;
      10'h167 : microOutput = 17'b00000000000000000;
      10'h168 : microOutput = 17'b00000000000000000;
      10'h169 : microOutput = 17'b00000000000000000;
      10'h16a : microOutput = 17'b00000000000000000;
      10'h16b : microOutput = 17'b00000000000000000;
      10'h16c : microOutput = 17'b00000000000000000;
      10'h16d : microOutput = 17'b00000000000000000;
      10'h16e : microOutput = 17'b00000000000000000;
      10'h16f : microOutput = 17'b00000000000000000;
      10'h170 : microOutput = 17'b10000000000000100;
      10'h171 : microOutput = 17'b00000000000000100;
      10'h172 : microOutput = 17'b00000100111000000;
      10'h173 : microOutput = 17'b00000100111000000;
      10'h174 : microOutput = 17'b00000100111000000;
      10'h175 : microOutput = 17'b00001100010101010;
      10'h176 : microOutput = 17'b00001000000010110;
      10'h177 : microOutput = 17'b00101001010000000;
      10'h178 : microOutput = 17'b10011000100000000;
      10'h179 : microOutput = 17'b00011011100100000;
      10'h17a : microOutput = 17'b01000100010000000;
      10'h17b : microOutput = 17'b01000000000001100;
      10'h17c : microOutput = 17'b10011000010000001;
      10'h17d : microOutput = 17'b10011011110100000;
      10'h17e : microOutput = 17'b10011111110100001;
      10'h17f : microOutput = 17'b00011000010000000;
      10'h180 : microOutput = 17'b00000000000000000;
      10'h181 : microOutput = 17'b00000000000000000;
      10'h182 : microOutput = 17'b00000000000000000;
      10'h183 : microOutput = 17'b00000000000000000;
      10'h184 : microOutput = 17'b00000000000000000;
      10'h185 : microOutput = 17'b00000000000000000;
      10'h186 : microOutput = 17'b00000000000000000;
      10'h187 : microOutput = 17'b00000000000000000;
      10'h188 : microOutput = 17'b00000000000000000;
      10'h189 : microOutput = 17'b00000000000000000;
      10'h18a : microOutput = 17'b00000000000000000;
      10'h18b : microOutput = 17'b00000000000000000;
      10'h18c : microOutput = 17'b00000000000000000;
      10'h18d : microOutput = 17'b00000000000000000;
      10'h18e : microOutput = 17'b00000000000000000;
      10'h18f : microOutput = 17'b00000000000000000;
      10'h190 : microOutput = 17'b00000000000000000;
      10'h191 : microOutput = 17'b00000000000000000;
      10'h192 : microOutput = 17'b00000000000000000;
      10'h193 : microOutput = 17'b00000000000000000;
      10'h194 : microOutput = 17'b00000000000000000;
      10'h195 : microOutput = 17'b00000000000000000;
      10'h196 : microOutput = 17'b00000000000000000;
      10'h197 : microOutput = 17'b00000000000000000;
      10'h198 : microOutput = 17'b00000000000000000;
      10'h199 : microOutput = 17'b00000000000000000;
      10'h19a : microOutput = 17'b00000000000000000;
      10'h19b : microOutput = 17'b00000000000000000;
      10'h19c : microOutput = 17'b00000000000000000;
      10'h19d : microOutput = 17'b00000000000000000;
      10'h19e : microOutput = 17'b00000000000000000;
      10'h19f : microOutput = 17'b00000000000000000;
      10'h1a0 : microOutput = 17'b00000000000000000;
      10'h1a1 : microOutput = 17'b00000000000000000;
      10'h1a2 : microOutput = 17'b00000000000000000;
      10'h1a3 : microOutput = 17'b00000000000000000;
      10'h1a4 : microOutput = 17'b00000000000000000;
      10'h1a5 : microOutput = 17'b00000000000000000;
      10'h1a6 : microOutput = 17'b00000000000000000;
      10'h1a7 : microOutput = 17'b00000000000000000;
      10'h1a8 : microOutput = 17'b00000000000000000;
      10'h1a9 : microOutput = 17'b00000000000000000;
      10'h1aa : microOutput = 17'b00000000000000000;
      10'h1ab : microOutput = 17'b00000000000000000;
      10'h1ac : microOutput = 17'b00000000000000000;
      10'h1ad : microOutput = 17'b00000000000000000;
      10'h1ae : microOutput = 17'b00000000000000000;
      10'h1af : microOutput = 17'b00000000000000000;
      10'h1b0 : microOutput = 17'b00000000000000000;
      10'h1b1 : microOutput = 17'b00000000000000000;
      10'h1b2 : microOutput = 17'b00000000000000000;
      10'h1b3 : microOutput = 17'b00000000000000000;
      10'h1b4 : microOutput = 17'b00000000000000000;
      10'h1b5 : microOutput = 17'b00000000000000000;
      10'h1b6 : microOutput = 17'b00000000000000000;
      10'h1b7 : microOutput = 17'b00000000000000000;
      10'h1b8 : microOutput = 17'b00000000000000000;
      10'h1b9 : microOutput = 17'b00000000000000000;
      10'h1ba : microOutput = 17'b00000000000000000;
      10'h1bb : microOutput = 17'b00000000000000000;
      10'h1bc : microOutput = 17'b00000000000000000;
      10'h1bd : microOutput = 17'b00000000000000000;
      10'h1be : microOutput = 17'b00000000000000000;
      10'h1bf : microOutput = 17'b00000000000000000;
      10'h1c0 : microOutput = 17'b00111110001000000;
      10'h1c1 : microOutput = 17'b10101011100100001;
      10'h1c2 : microOutput = 17'b10001010100000000;
      10'h1c3 : microOutput = 17'b10101011100100001;
      10'h1c4 : microOutput = 17'b00100011010000000;
      10'h1c5 : microOutput = 17'b10110000001100001;
      10'h1c6 : microOutput = 17'b10000000110000000;
      10'h1c7 : microOutput = 17'b10110000101100001;
      10'h1c8 : microOutput = 17'b00000000000000000;
      10'h1c9 : microOutput = 17'b10110000101100001;
      10'h1ca : microOutput = 17'b10110110110100000;
      10'h1cb : microOutput = 17'b10100001110100001;
      10'h1cc : microOutput = 17'b00111100010000000;
      10'h1cd : microOutput = 17'b10011101100000001;
      10'h1ce : microOutput = 17'b10111110100100000;
      10'h1cf : microOutput = 17'b10010011010100001;
      10'h1d0 : microOutput = 17'b00111100010100000;
      10'h1d1 : microOutput = 17'b10101011100000001;
      10'h1d2 : microOutput = 17'b10101001101000000;
      10'h1d3 : microOutput = 17'b10101011100000001;
      10'h1d4 : microOutput = 17'b00000000000000000;
      10'h1d5 : microOutput = 17'b10011111000100001;
      10'h1d6 : microOutput = 17'b10101001111000000;
      10'h1d7 : microOutput = 17'b10011011000100001;
      10'h1d8 : microOutput = 17'b00000000000000000;
      10'h1d9 : microOutput = 17'b10010011010100001;
      10'h1da : microOutput = 17'b00000000000000000;
      10'h1db : microOutput = 17'b00000000000000000;
      10'h1dc : microOutput = 17'b00000000000000000;
      10'h1dd : microOutput = 17'b00000000000000000;
      10'h1de : microOutput = 17'b00000000000000000;
      10'h1df : microOutput = 17'b00000000000000000;
      10'h1e0 : microOutput = 17'b00001010100000000;
      10'h1e1 : microOutput = 17'b10111110000100000;
      10'h1e2 : microOutput = 17'b10000100100000000;
      10'h1e3 : microOutput = 17'b00111010001100000;
      10'h1e4 : microOutput = 17'b00000000110000000;
      10'h1e5 : microOutput = 17'b10011001000000000;
      10'h1e6 : microOutput = 17'b10000100110000000;
      10'h1e7 : microOutput = 17'b00111010011100000;
      10'h1e8 : microOutput = 17'b00101101101100000;
      10'h1e9 : microOutput = 17'b10001110111000000;
      10'h1ea : microOutput = 17'b10101111101000000;
      10'h1eb : microOutput = 17'b00010100100000000;
      10'h1ec : microOutput = 17'b00101011111000000;
      10'h1ed : microOutput = 17'b10110100001100000;
      10'h1ee : microOutput = 17'b10101111111000000;
      10'h1ef : microOutput = 17'b00010100010000000;
      10'h1f0 : microOutput = 17'b00111000100000000;
      10'h1f1 : microOutput = 17'b10110100101100000;
      10'h1f2 : microOutput = 17'b10101001010100000;
      10'h1f3 : microOutput = 17'b00101011001000000;
      10'h1f4 : microOutput = 17'b00100001100000000;
      10'h1f5 : microOutput = 17'b10001110010000000;
      10'h1f6 : microOutput = 17'b10101111001000000;
      10'h1f7 : microOutput = 17'b00101011011000000;
      10'h1f8 : microOutput = 17'b00000110010111010;
      10'h1f9 : microOutput = 17'b10111000110000000;
      10'h1fa : microOutput = 17'b10011101110100000;
      10'h1fb : microOutput = 17'b00111010101100000;
      10'h1fc : microOutput = 17'b00000000000000000;
      10'h1fd : microOutput = 17'b10101011011100000;
      10'h1fe : microOutput = 17'b01100011110100001;
      10'h1ff : microOutput = 17'b00111010111100000;
      10'h200 : microOutput = 17'b00000000000000000;
      10'h201 : microOutput = 17'b00000000000000000;
      10'h202 : microOutput = 17'b00000000000000000;
      10'h203 : microOutput = 17'b00000000000000000;
      10'h204 : microOutput = 17'b00000000000000000;
      10'h205 : microOutput = 17'b00000000000000000;
      10'h206 : microOutput = 17'b00000000000000000;
      10'h207 : microOutput = 17'b00000000000000000;
      10'h208 : microOutput = 17'b00000000000000000;
      10'h209 : microOutput = 17'b00000000000000000;
      10'h20a : microOutput = 17'b00000000000000000;
      10'h20b : microOutput = 17'b00000000000000000;
      10'h20c : microOutput = 17'b00000000000000000;
      10'h20d : microOutput = 17'b00000000000000000;
      10'h20e : microOutput = 17'b00000000000000000;
      10'h20f : microOutput = 17'b00000000000000000;
      10'h210 : microOutput = 17'b00100101000000000;
      10'h211 : microOutput = 17'b00000100000010110;
      10'h212 : microOutput = 17'b00000000000000100;
      10'h213 : microOutput = 17'b00001110000001110;
      10'h214 : microOutput = 17'b00100001000000000;
      10'h215 : microOutput = 17'b10110000110100001;
      10'h216 : microOutput = 17'b00100101011001010;
      10'h217 : microOutput = 17'b00111000001100000;
      10'h218 : microOutput = 17'b00100101100000001;
      10'h219 : microOutput = 17'b10011000010000000;
      10'h21a : microOutput = 17'b01101101100000000;
      10'h21b : microOutput = 17'b00000000000001100;
      10'h21c : microOutput = 17'b01100101110000000;
      10'h21d : microOutput = 17'b00000000000001100;
      10'h21e : microOutput = 17'b00001100001111010;
      10'h21f : microOutput = 17'b01001100001111010;
      10'h220 : microOutput = 17'b00000000000000000;
      10'h221 : microOutput = 17'b00000000000000000;
      10'h222 : microOutput = 17'b00000000000000000;
      10'h223 : microOutput = 17'b00000000000000000;
      10'h224 : microOutput = 17'b00000000000000000;
      10'h225 : microOutput = 17'b00000000000000000;
      10'h226 : microOutput = 17'b00000000000000000;
      10'h227 : microOutput = 17'b00000000000000000;
      10'h228 : microOutput = 17'b00000000000000000;
      10'h229 : microOutput = 17'b00000000000000000;
      10'h22a : microOutput = 17'b00000000000000000;
      10'h22b : microOutput = 17'b00000000000000000;
      10'h22c : microOutput = 17'b00000000000000000;
      10'h22d : microOutput = 17'b00000000000000000;
      10'h22e : microOutput = 17'b00000000000000000;
      10'h22f : microOutput = 17'b00000000000000000;
      10'h230 : microOutput = 17'b10101111000000001;
      10'h231 : microOutput = 17'b00000100111000000;
      10'h232 : microOutput = 17'b10101111000000001;
      10'h233 : microOutput = 17'b00000000000000100;
      10'h234 : microOutput = 17'b00100111010000000;
      10'h235 : microOutput = 17'b00001110101100000;
      10'h236 : microOutput = 17'b11010001100000000;
      10'h237 : microOutput = 17'b00110010100111010;
      10'h238 : microOutput = 17'b00000000000000100;
      10'h239 : microOutput = 17'b00000100111000000;
      10'h23a : microOutput = 17'b00000000000000100;
      10'h23b : microOutput = 17'b10110000110100001;
      10'h23c : microOutput = 17'b01100111110000001;
      10'h23d : microOutput = 17'b10000000000000100;
      10'h23e : microOutput = 17'b01111100100100000;
      10'h23f : microOutput = 17'b01100001100100001;
      10'h240 : microOutput = 17'b00000000000000000;
      10'h241 : microOutput = 17'b00000000000000000;
      10'h242 : microOutput = 17'b00000000000000000;
      10'h243 : microOutput = 17'b00000000000000000;
      10'h244 : microOutput = 17'b00000000000000000;
      10'h245 : microOutput = 17'b00000000000000000;
      10'h246 : microOutput = 17'b00000000000000000;
      10'h247 : microOutput = 17'b00000000000000000;
      10'h248 : microOutput = 17'b00000000000000000;
      10'h249 : microOutput = 17'b00000000000000000;
      10'h24a : microOutput = 17'b00000000000000000;
      10'h24b : microOutput = 17'b00000000000000000;
      10'h24c : microOutput = 17'b00000000000000000;
      10'h24d : microOutput = 17'b00000000000000000;
      10'h24e : microOutput = 17'b00000000000000000;
      10'h24f : microOutput = 17'b00000000000000000;
      10'h250 : microOutput = 17'b00000000001100000;
      10'h251 : microOutput = 17'b10001010010100001;
      10'h252 : microOutput = 17'b00110110100000110;
      10'h253 : microOutput = 17'b00000000000000100;
      10'h254 : microOutput = 17'b00100001000000000;
      10'h255 : microOutput = 17'b10111110000100000;
      10'h256 : microOutput = 17'b10100111000100000;
      10'h257 : microOutput = 17'b00111000010000000;
      10'h258 : microOutput = 17'b10000000000000100;
      10'h259 : microOutput = 17'b00101001100100000;
      10'h25a : microOutput = 17'b00101101100100000;
      10'h25b : microOutput = 17'b00000000000000100;
      10'h25c : microOutput = 17'b00100101110100000;
      10'h25d : microOutput = 17'b00000000000000100;
      10'h25e : microOutput = 17'b00100101110100000;
      10'h25f : microOutput = 17'b00100101110100000;
      10'h260 : microOutput = 17'b00000000000000000;
      10'h261 : microOutput = 17'b00000000000000000;
      10'h262 : microOutput = 17'b00000000000000000;
      10'h263 : microOutput = 17'b00000000000000000;
      10'h264 : microOutput = 17'b00000000000000000;
      10'h265 : microOutput = 17'b00000000000000000;
      10'h266 : microOutput = 17'b00000000000000000;
      10'h267 : microOutput = 17'b00000000000000000;
      10'h268 : microOutput = 17'b00000000000000000;
      10'h269 : microOutput = 17'b00000000000000000;
      10'h26a : microOutput = 17'b00000000000000000;
      10'h26b : microOutput = 17'b00000000000000000;
      10'h26c : microOutput = 17'b00000000000000000;
      10'h26d : microOutput = 17'b00000000000000000;
      10'h26e : microOutput = 17'b00000000000000000;
      10'h26f : microOutput = 17'b00000000000000000;
      10'h270 : microOutput = 17'b10100111000100000;
      10'h271 : microOutput = 17'b01101011000100000;
      10'h272 : microOutput = 17'b01111110000100001;
      10'h273 : microOutput = 17'b10100111000100000;
      10'h274 : microOutput = 17'b10100111001000000;
      10'h275 : microOutput = 17'b10111110000100000;
      10'h276 : microOutput = 17'b00101111010000000;
      10'h277 : microOutput = 17'b00110010100111010;
      10'h278 : microOutput = 17'b00000000000000100;
      10'h279 : microOutput = 17'b10100011100100001;
      10'h27a : microOutput = 17'b00000000000000100;
      10'h27b : microOutput = 17'b00000010011100001;
      10'h27c : microOutput = 17'b10100111110100000;
      10'h27d : microOutput = 17'b00000000000000100;
      10'h27e : microOutput = 17'b00101111110100000;
      10'h27f : microOutput = 17'b00101111101100000;
      10'h280 : microOutput = 17'b00000000000000000;
      10'h281 : microOutput = 17'b00000000000000000;
      10'h282 : microOutput = 17'b00000000000000000;
      10'h283 : microOutput = 17'b00000000000000000;
      10'h284 : microOutput = 17'b00000000000000000;
      10'h285 : microOutput = 17'b00000000000000000;
      10'h286 : microOutput = 17'b00000000000000000;
      10'h287 : microOutput = 17'b00000000000000000;
      10'h288 : microOutput = 17'b00000000000000000;
      10'h289 : microOutput = 17'b00000000000000000;
      10'h28a : microOutput = 17'b00000000000000000;
      10'h28b : microOutput = 17'b00000000000000000;
      10'h28c : microOutput = 17'b00000000000000000;
      10'h28d : microOutput = 17'b00000000000000000;
      10'h28e : microOutput = 17'b00000000000000000;
      10'h28f : microOutput = 17'b00000000000000000;
      10'h290 : microOutput = 17'b00100101001000000;
      10'h291 : microOutput = 17'b00101001000010110;
      10'h292 : microOutput = 17'b00110010000100000;
      10'h293 : microOutput = 17'b00100011000100000;
      10'h294 : microOutput = 17'b00100101011000000;
      10'h295 : microOutput = 17'b00101001011100000;
      10'h296 : microOutput = 17'b00101011110110000;
      10'h297 : microOutput = 17'b00101111001000000;
      10'h298 : microOutput = 17'b00010100000000000;
      10'h299 : microOutput = 17'b10110100111000001;
      10'h29a : microOutput = 17'b01110010100100000;
      10'h29b : microOutput = 17'b10110000110100001;
      10'h29c : microOutput = 17'b00010100110000000;
      10'h29d : microOutput = 17'b10110100110100001;
      10'h29e : microOutput = 17'b01111000110100000;
      10'h29f : microOutput = 17'b10111110110100001;
      10'h2a0 : microOutput = 17'b00000000000000000;
      10'h2a1 : microOutput = 17'b00000000000000000;
      10'h2a2 : microOutput = 17'b00000000000000000;
      10'h2a3 : microOutput = 17'b00000000000000000;
      10'h2a4 : microOutput = 17'b00000000000000000;
      10'h2a5 : microOutput = 17'b00000000000000000;
      10'h2a6 : microOutput = 17'b00000000000000000;
      10'h2a7 : microOutput = 17'b00000000000000000;
      10'h2a8 : microOutput = 17'b00000000000000000;
      10'h2a9 : microOutput = 17'b00000000000000000;
      10'h2aa : microOutput = 17'b00000000000000000;
      10'h2ab : microOutput = 17'b00000000000000000;
      10'h2ac : microOutput = 17'b00000000000000000;
      10'h2ad : microOutput = 17'b00000000000000000;
      10'h2ae : microOutput = 17'b00000000000000000;
      10'h2af : microOutput = 17'b00000000000000000;
      10'h2b0 : microOutput = 17'b00100011010100000;
      10'h2b1 : microOutput = 17'b00100111000100000;
      10'h2b2 : microOutput = 17'b00000110100000010;
      10'h2b3 : microOutput = 17'b10111110000100000;
      10'h2b4 : microOutput = 17'b00000100011100000;
      10'h2b5 : microOutput = 17'b00110000110000000;
      10'h2b6 : microOutput = 17'b00000110110000010;
      10'h2b7 : microOutput = 17'b10010001110000000;
      10'h2b8 : microOutput = 17'b10110100111000001;
      10'h2b9 : microOutput = 17'b10000000000001000;
      10'h2ba : microOutput = 17'b01110000100100000;
      10'h2bb : microOutput = 17'b10110100101000000;
      10'h2bc : microOutput = 17'b10010101110100001;
      10'h2bd : microOutput = 17'b10111110000100000;
      10'h2be : microOutput = 17'b01101101111100000;
      10'h2bf : microOutput = 17'b10101011101000000;
      10'h2c0 : microOutput = 17'b00000000000000000;
      10'h2c1 : microOutput = 17'b00000000000000000;
      10'h2c2 : microOutput = 17'b00000000000000000;
      10'h2c3 : microOutput = 17'b00000000000000000;
      10'h2c4 : microOutput = 17'b00000000000000000;
      10'h2c5 : microOutput = 17'b00000000000000000;
      10'h2c6 : microOutput = 17'b00000000000000000;
      10'h2c7 : microOutput = 17'b00000000000000000;
      10'h2c8 : microOutput = 17'b00000000000000000;
      10'h2c9 : microOutput = 17'b00000000000000000;
      10'h2ca : microOutput = 17'b00000000000000000;
      10'h2cb : microOutput = 17'b00000000000000000;
      10'h2cc : microOutput = 17'b00000000000000000;
      10'h2cd : microOutput = 17'b00000000000000000;
      10'h2ce : microOutput = 17'b00000000000000000;
      10'h2cf : microOutput = 17'b00000000000000000;
      10'h2d0 : microOutput = 17'b00101001000010110;
      10'h2d1 : microOutput = 17'b10001010011100001;
      10'h2d2 : microOutput = 17'b00100001000000110;
      10'h2d3 : microOutput = 17'b00101101000000110;
      10'h2d4 : microOutput = 17'b00101001011100000;
      10'h2d5 : microOutput = 17'b10001010011100001;
      10'h2d6 : microOutput = 17'b00110110111000110;
      10'h2d7 : microOutput = 17'b00101101010000110;
      10'h2d8 : microOutput = 17'b10001100101000001;
      10'h2d9 : microOutput = 17'b10110100101000000;
      10'h2da : microOutput = 17'b10101101101100000;
      10'h2db : microOutput = 17'b01111110000100001;
      10'h2dc : microOutput = 17'b10100101100100001;
      10'h2dd : microOutput = 17'b10101011101000000;
      10'h2de : microOutput = 17'b10101011111000000;
      10'h2df : microOutput = 17'b01100001100100001;
      10'h2e0 : microOutput = 17'b00000000000000000;
      10'h2e1 : microOutput = 17'b00000000000000000;
      10'h2e2 : microOutput = 17'b00000000000000000;
      10'h2e3 : microOutput = 17'b00000000000000000;
      10'h2e4 : microOutput = 17'b00000000000000000;
      10'h2e5 : microOutput = 17'b00000000000000000;
      10'h2e6 : microOutput = 17'b00000000000000000;
      10'h2e7 : microOutput = 17'b00000000000000000;
      10'h2e8 : microOutput = 17'b00000000000000000;
      10'h2e9 : microOutput = 17'b00000000000000000;
      10'h2ea : microOutput = 17'b00000000000000000;
      10'h2eb : microOutput = 17'b00000000000000000;
      10'h2ec : microOutput = 17'b00000000000000000;
      10'h2ed : microOutput = 17'b00000000000000000;
      10'h2ee : microOutput = 17'b00000000000000000;
      10'h2ef : microOutput = 17'b00000000000000000;
      10'h2f0 : microOutput = 17'b00110010100111010;
      10'h2f1 : microOutput = 17'b10001010010100001;
      10'h2f2 : microOutput = 17'b10110100100000000;
      10'h2f3 : microOutput = 17'b10110100111000001;
      10'h2f4 : microOutput = 17'b01110010110111010;
      10'h2f5 : microOutput = 17'b10001010010100001;
      10'h2f6 : microOutput = 17'b10101011010100000;
      10'h2f7 : microOutput = 17'b10110100110100001;
      10'h2f8 : microOutput = 17'b10111100100100001;
      10'h2f9 : microOutput = 17'b01101111110000000;
      10'h2fa : microOutput = 17'b01000110010000001;
      10'h2fb : microOutput = 17'b10101111111100000;
      10'h2fc : microOutput = 17'b10101011110000001;
      10'h2fd : microOutput = 17'b01100011110000000;
      10'h2fe : microOutput = 17'b01110100100100001;
      10'h2ff : microOutput = 17'b10110000000000000;
      10'h300 : microOutput = 17'b10011001110000000;
      10'h301 : microOutput = 17'b00110110000000000;
      10'h302 : microOutput = 17'b00101111001000000;
      10'h303 : microOutput = 17'b10111110000100000;
      10'h304 : microOutput = 17'b00110100111000000;
      10'h305 : microOutput = 17'b10001100100100000;
      10'h306 : microOutput = 17'b00000000000000100;
      10'h307 : microOutput = 17'b00110010000000000;
      10'h308 : microOutput = 17'b00000100010100110;
      10'h309 : microOutput = 17'b00111110000100000;
      10'h30a : microOutput = 17'b00111110000100000;
      10'h30b : microOutput = 17'b10100111011000000;
      10'h30c : microOutput = 17'b01110100110000001;
      10'h30d : microOutput = 17'b01110100100100000;
      10'h30e : microOutput = 17'b10010101000000000;
      10'h30f : microOutput = 17'b10110110100000000;
      10'h310 : microOutput = 17'b00000000000000000;
      10'h311 : microOutput = 17'b00000000000000000;
      10'h312 : microOutput = 17'b00000000000000000;
      10'h313 : microOutput = 17'b00000000000000000;
      10'h314 : microOutput = 17'b00000000000000000;
      10'h315 : microOutput = 17'b00000000000000000;
      10'h316 : microOutput = 17'b00000000000000000;
      10'h317 : microOutput = 17'b00000000000000000;
      10'h318 : microOutput = 17'b00000000000000000;
      10'h319 : microOutput = 17'b00000000000000000;
      10'h31a : microOutput = 17'b00000000000000000;
      10'h31b : microOutput = 17'b00000000000000000;
      10'h31c : microOutput = 17'b00000000000000000;
      10'h31d : microOutput = 17'b00000000000000000;
      10'h31e : microOutput = 17'b00000000000000000;
      10'h31f : microOutput = 17'b00000000000000000;
      10'h320 : microOutput = 17'b00110110000000000;
      10'h321 : microOutput = 17'b00010110001100000;
      10'h322 : microOutput = 17'b00000110010111010;
      10'h323 : microOutput = 17'b00000110010111010;
      10'h324 : microOutput = 17'b00110100111000000;
      10'h325 : microOutput = 17'b10111010010000000;
      10'h326 : microOutput = 17'b00001110110000000;
      10'h327 : microOutput = 17'b00000000000000100;
      10'h328 : microOutput = 17'b10110000110100001;
      10'h329 : microOutput = 17'b01111010100000000;
      10'h32a : microOutput = 17'b01010110001100001;
      10'h32b : microOutput = 17'b10111010110000000;
      10'h32c : microOutput = 17'b10110000110100000;
      10'h32d : microOutput = 17'b00100001010001010;
      10'h32e : microOutput = 17'b01010110001100001;
      10'h32f : microOutput = 17'b01110000100100000;
      10'h330 : microOutput = 17'b00000000000000000;
      10'h331 : microOutput = 17'b00000000000000000;
      10'h332 : microOutput = 17'b00000000000000000;
      10'h333 : microOutput = 17'b00000000000000000;
      10'h334 : microOutput = 17'b00000000000000000;
      10'h335 : microOutput = 17'b00000000000000000;
      10'h336 : microOutput = 17'b00000000000000000;
      10'h337 : microOutput = 17'b00000000000000000;
      10'h338 : microOutput = 17'b00000000000000000;
      10'h339 : microOutput = 17'b00000000000000000;
      10'h33a : microOutput = 17'b00000000000000000;
      10'h33b : microOutput = 17'b00000000000000000;
      10'h33c : microOutput = 17'b00000000000000000;
      10'h33d : microOutput = 17'b00000000000000000;
      10'h33e : microOutput = 17'b00000000000000000;
      10'h33f : microOutput = 17'b00000000000000000;
      10'h340 : microOutput = 17'b00000100111000000;
      10'h341 : microOutput = 17'b10111000000100001;
      10'h342 : microOutput = 17'b00000000000000100;
      10'h343 : microOutput = 17'b00110000010100000;
      10'h344 : microOutput = 17'b01111110000100000;
      10'h345 : microOutput = 17'b10111000010100001;
      10'h346 : microOutput = 17'b00000000000000100;
      10'h347 : microOutput = 17'b00111000001100000;
      10'h348 : microOutput = 17'b01111110000100000;
      10'h349 : microOutput = 17'b10000000000000100;
      10'h34a : microOutput = 17'b01111100100100000;
      10'h34b : microOutput = 17'b01000000000000100;
      10'h34c : microOutput = 17'b00000000000000100;
      10'h34d : microOutput = 17'b01110100111000000;
      10'h34e : microOutput = 17'b01111100110100000;
      10'h34f : microOutput = 17'b01110010100100000;
      10'h350 : microOutput = 17'b00000000000000000;
      10'h351 : microOutput = 17'b00000000000000000;
      10'h352 : microOutput = 17'b00000000000000000;
      10'h353 : microOutput = 17'b00000000000000000;
      10'h354 : microOutput = 17'b00000000000000000;
      10'h355 : microOutput = 17'b00000000000000000;
      10'h356 : microOutput = 17'b00000000000000000;
      10'h357 : microOutput = 17'b00000000000000000;
      10'h358 : microOutput = 17'b00000000000000000;
      10'h359 : microOutput = 17'b00000000000000000;
      10'h35a : microOutput = 17'b00000000000000000;
      10'h35b : microOutput = 17'b00000000000000000;
      10'h35c : microOutput = 17'b00000000000000000;
      10'h35d : microOutput = 17'b00000000000000000;
      10'h35e : microOutput = 17'b00000000000000000;
      10'h35f : microOutput = 17'b00000000000000000;
      10'h360 : microOutput = 17'b01001110111100000;
      10'h361 : microOutput = 17'b00000000000000100;
      10'h362 : microOutput = 17'b00000000000000100;
      10'h363 : microOutput = 17'b10110000110100001;
      10'h364 : microOutput = 17'b00000000000000000;
      10'h365 : microOutput = 17'b00000000000000000;
      10'h366 : microOutput = 17'b00000000000000000;
      10'h367 : microOutput = 17'b01011001100000000;
      10'h368 : microOutput = 17'b01111010100100001;
      10'h369 : microOutput = 17'b00000000001001010;
      10'h36a : microOutput = 17'b10000000000000100;
      10'h36b : microOutput = 17'b01110010110100000;
      10'h36c : microOutput = 17'b01110110110100000;
      10'h36d : microOutput = 17'b01111010110100001;
      10'h36e : microOutput = 17'b01111110000100000;
      10'h36f : microOutput = 17'b00000000000000100;
      10'h370 : microOutput = 17'b00000000000000000;
      10'h371 : microOutput = 17'b00000000000000000;
      10'h372 : microOutput = 17'b00000000000000000;
      10'h373 : microOutput = 17'b00000000000000000;
      10'h374 : microOutput = 17'b00000000000000000;
      10'h375 : microOutput = 17'b00000000000000000;
      10'h376 : microOutput = 17'b00000000000000000;
      10'h377 : microOutput = 17'b00000000000000000;
      10'h378 : microOutput = 17'b00000000000000000;
      10'h379 : microOutput = 17'b00000000000000000;
      10'h37a : microOutput = 17'b00000000000000000;
      10'h37b : microOutput = 17'b00000000000000000;
      10'h37c : microOutput = 17'b00000000000000000;
      10'h37d : microOutput = 17'b00000000000000000;
      10'h37e : microOutput = 17'b00000000000000000;
      10'h37f : microOutput = 17'b00000000000000000;
      10'h380 : microOutput = 17'b10001100110100111;
      10'h381 : microOutput = 17'b10111100001000001;
      10'h382 : microOutput = 17'b10111100001000001;
      10'h383 : microOutput = 17'b00101101000000110;
      10'h384 : microOutput = 17'b10001100101100111;
      10'h385 : microOutput = 17'b10111100011000001;
      10'h386 : microOutput = 17'b10111100011000001;
      10'h387 : microOutput = 17'b00101101010000110;
      10'h388 : microOutput = 17'b10110100101000000;
      10'h389 : microOutput = 17'b01111110000100000;
      10'h38a : microOutput = 17'b10110100101000000;
      10'h38b : microOutput = 17'b10111100100100001;
      10'h38c : microOutput = 17'b10111110110000000;
      10'h38d : microOutput = 17'b01000000000000100;
      10'h38e : microOutput = 17'b10111110110000000;
      10'h38f : microOutput = 17'b10111000100100001;
      10'h390 : microOutput = 17'b00000000000000000;
      10'h391 : microOutput = 17'b00000000000000000;
      10'h392 : microOutput = 17'b00000000000000000;
      10'h393 : microOutput = 17'b00000000000000000;
      10'h394 : microOutput = 17'b00000000000000000;
      10'h395 : microOutput = 17'b00000000000000000;
      10'h396 : microOutput = 17'b00000000000000000;
      10'h397 : microOutput = 17'b00000000000000000;
      10'h398 : microOutput = 17'b00000000000000000;
      10'h399 : microOutput = 17'b00000000000000000;
      10'h39a : microOutput = 17'b00000000000000000;
      10'h39b : microOutput = 17'b00000000000000000;
      10'h39c : microOutput = 17'b00000000000000000;
      10'h39d : microOutput = 17'b00000000000000000;
      10'h39e : microOutput = 17'b00000000000000000;
      10'h39f : microOutput = 17'b00000000000000000;
      10'h3a0 : microOutput = 17'b10111110000000000;
      10'h3a1 : microOutput = 17'b10110010010000001;
      10'h3a2 : microOutput = 17'b00111110010000001;
      10'h3a3 : microOutput = 17'b00111000001100000;
      10'h3a4 : microOutput = 17'b10101001110000000;
      10'h3a5 : microOutput = 17'b10110000000100001;
      10'h3a6 : microOutput = 17'b00101111100100000;
      10'h3a7 : microOutput = 17'b00111000101110000;
      10'h3a8 : microOutput = 17'b00110010100111010;
      10'h3a9 : microOutput = 17'b01111010101000000;
      10'h3aa : microOutput = 17'b01000110010000001;
      10'h3ab : microOutput = 17'b01000110010000000;
      10'h3ac : microOutput = 17'b01110010110111010;
      10'h3ad : microOutput = 17'b01111010111000000;
      10'h3ae : microOutput = 17'b01110100100100001;
      10'h3af : microOutput = 17'b01110100100100001;
      10'h3b0 : microOutput = 17'b00000000000000000;
      10'h3b1 : microOutput = 17'b00000000000000000;
      10'h3b2 : microOutput = 17'b00000000000000000;
      10'h3b3 : microOutput = 17'b00000000000000000;
      10'h3b4 : microOutput = 17'b00000000000000000;
      10'h3b5 : microOutput = 17'b00000000000000000;
      10'h3b6 : microOutput = 17'b00000000000000000;
      10'h3b7 : microOutput = 17'b00000000000000000;
      10'h3b8 : microOutput = 17'b00000000000000000;
      10'h3b9 : microOutput = 17'b00000000000000000;
      10'h3ba : microOutput = 17'b00000000000000000;
      10'h3bb : microOutput = 17'b00000000000000000;
      10'h3bc : microOutput = 17'b00000000000000000;
      10'h3bd : microOutput = 17'b00000000000000000;
      10'h3be : microOutput = 17'b00000000000000000;
      10'h3bf : microOutput = 17'b00000000000000000;
      10'h3c0 : microOutput = 17'b00101001110100000;
      10'h3c1 : microOutput = 17'b10001100100100000;
      10'h3c2 : microOutput = 17'b01110010000100000;
      10'h3c3 : microOutput = 17'b10110000110100001;
      10'h3c4 : microOutput = 17'b00000010000011110;
      10'h3c5 : microOutput = 17'b01111000000000000;
      10'h3c6 : microOutput = 17'b01000000101000000;
      10'h3c7 : microOutput = 17'b10110000010000001;
      10'h3c8 : microOutput = 17'b00101101110100000;
      10'h3c9 : microOutput = 17'b10111010000000000;
      10'h3ca : microOutput = 17'b01001010001000000;
      10'h3cb : microOutput = 17'b10110110000100001;
      10'h3cc : microOutput = 17'b00000000000000000;
      10'h3cd : microOutput = 17'b00000000000000000;
      10'h3ce : microOutput = 17'b00000000000000000;
      10'h3cf : microOutput = 17'b00000000000000000;
      10'h3d0 : microOutput = 17'b00000000000000000;
      10'h3d1 : microOutput = 17'b00000000000000000;
      10'h3d2 : microOutput = 17'b00000000000000000;
      10'h3d3 : microOutput = 17'b00000000000000000;
      10'h3d4 : microOutput = 17'b00000000000000000;
      10'h3d5 : microOutput = 17'b00000000000000000;
      10'h3d6 : microOutput = 17'b00000000000000000;
      10'h3d7 : microOutput = 17'b00000000000000000;
      10'h3d8 : microOutput = 17'b00000000000000000;
      10'h3d9 : microOutput = 17'b00000000000000000;
      10'h3da : microOutput = 17'b00000000000000000;
      10'h3db : microOutput = 17'b00000000000000000;
      10'h3dc : microOutput = 17'b00000000000000000;
      10'h3dd : microOutput = 17'b00000000000000000;
      10'h3de : microOutput = 17'b00000000000000000;
      10'h3df : microOutput = 17'b00000000000000000;
      10'h3e0 : microOutput = 17'b10100111101000000;
      10'h3e1 : microOutput = 17'b00000000000000000;
      10'h3e2 : microOutput = 17'b10010010000000010;
      10'h3e3 : microOutput = 17'b10100111000000001;
      10'h3e4 : microOutput = 17'b10100111111000000;
      10'h3e5 : microOutput = 17'b00000000000000000;
      10'h3e6 : microOutput = 17'b10010010010000010;
      10'h3e7 : microOutput = 17'b10001110011100001;
      10'h3e8 : microOutput = 17'b00100011001100000;
      10'h3e9 : microOutput = 17'b00100001001001010;
      10'h3ea : microOutput = 17'b10010011000000010;
      10'h3eb : microOutput = 17'b10001010110100001;
      10'h3ec : microOutput = 17'b01100011011100000;
      10'h3ed : microOutput = 17'b00100001011001010;
      10'h3ee : microOutput = 17'b10010011010000010;
      10'h3ef : microOutput = 17'b10001010100100001;
      10'h3f0 : microOutput = 17'b00000000000000000;
      10'h3f1 : microOutput = 17'b00000000000000000;
      10'h3f2 : microOutput = 17'b00000000000000000;
      10'h3f3 : microOutput = 17'b00000000000000000;
      10'h3f4 : microOutput = 17'b00000000000000000;
      10'h3f5 : microOutput = 17'b00000000000000000;
      10'h3f6 : microOutput = 17'b00000000000000000;
      10'h3f7 : microOutput = 17'b00000000000000000;
      10'h3f8 : microOutput = 17'b00000000000000000;
      10'h3f9 : microOutput = 17'b00000000000000000;
      10'h3fa : microOutput = 17'b00000000000000000;
      10'h3fb : microOutput = 17'b00000000000000000;
      10'h3fc : microOutput = 17'b00000000000000000;
      10'h3fd : microOutput = 17'b00000000000000000;
      10'h3fe : microOutput = 17'b00000000000000000;
      10'h3ff : microOutput = 17'b00000000000000000;
      default : ;
    endcase
  end

endmodule
